VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO skullart
  CLASS BLOCK ;
  FOREIGN skullart ;
  ORIGIN -10.000 -10.000 ;
  SIZE 140.000 BY 160.000 ;
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 10.000 10.000 15.000 170.000 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 145.000 10.000 150.000 170.000 ;
    END
  END vccd1
  OBS
      LAYER met1 ;
        RECT 83.000 164.000 84.000 165.000 ;
        RECT 93.000 164.000 94.000 165.000 ;
        RECT 114.000 164.000 115.000 165.000 ;
        RECT 40.000 163.000 45.000 164.000 ;
        RECT 39.000 162.000 44.000 163.000 ;
        RECT 37.000 154.000 38.000 155.000 ;
        RECT 37.000 153.000 39.000 154.000 ;
        RECT 41.000 153.000 44.000 162.000 ;
        RECT 49.000 162.000 59.000 164.000 ;
        RECT 49.000 160.000 52.000 162.000 ;
        RECT 50.000 159.000 52.000 160.000 ;
        RECT 51.000 158.000 52.000 159.000 ;
        RECT 56.000 157.000 59.000 162.000 ;
        RECT 69.000 157.000 72.000 164.000 ;
        RECT 75.000 163.000 84.000 164.000 ;
        RECT 75.000 162.000 77.000 163.000 ;
        RECT 79.000 162.000 84.000 163.000 ;
        RECT 75.000 161.000 76.000 162.000 ;
        RECT 53.000 156.000 61.000 157.000 ;
        RECT 66.000 156.000 74.000 157.000 ;
        RECT 53.000 155.000 60.000 156.000 ;
        RECT 66.000 155.000 73.000 156.000 ;
        RECT 51.000 153.000 52.000 154.000 ;
        RECT 37.000 152.000 45.000 153.000 ;
        RECT 50.000 152.000 52.000 153.000 ;
        RECT 37.000 151.000 47.000 152.000 ;
        RECT 38.000 150.000 48.000 151.000 ;
        RECT 49.000 150.000 52.000 152.000 ;
        RECT 56.000 150.000 59.000 155.000 ;
        RECT 64.000 153.000 65.000 154.000 ;
        RECT 63.000 152.000 65.000 153.000 ;
        RECT 62.000 150.000 65.000 152.000 ;
        RECT 69.000 150.000 72.000 155.000 ;
        RECT 81.000 150.000 84.000 162.000 ;
        RECT 85.000 163.000 94.000 164.000 ;
        RECT 97.000 163.000 105.000 164.000 ;
        RECT 107.000 163.000 108.000 164.000 ;
        RECT 85.000 162.000 87.000 163.000 ;
        RECT 89.000 162.000 94.000 163.000 ;
        RECT 96.000 162.000 105.000 163.000 ;
        RECT 85.000 161.000 86.000 162.000 ;
        RECT 91.000 150.000 94.000 162.000 ;
        RECT 95.000 150.000 98.000 162.000 ;
        RECT 41.000 148.000 44.000 150.000 ;
        RECT 49.000 149.000 58.000 150.000 ;
        RECT 62.000 149.000 71.000 150.000 ;
        RECT 81.000 149.000 83.000 150.000 ;
        RECT 91.000 149.000 93.000 150.000 ;
        RECT 96.000 149.000 98.000 150.000 ;
        RECT 49.000 148.000 57.000 149.000 ;
        RECT 62.000 148.000 70.000 149.000 ;
        RECT 81.000 148.000 82.000 149.000 ;
        RECT 91.000 148.000 92.000 149.000 ;
        RECT 97.000 148.000 98.000 149.000 ;
        RECT 102.000 148.000 105.000 162.000 ;
        RECT 106.000 162.000 109.000 163.000 ;
        RECT 106.000 161.000 110.000 162.000 ;
        RECT 107.000 160.000 111.000 161.000 ;
        RECT 108.000 159.000 111.000 160.000 ;
        RECT 109.000 158.000 111.000 159.000 ;
        RECT 112.000 158.000 115.000 164.000 ;
        RECT 120.000 163.000 129.000 164.000 ;
        RECT 119.000 162.000 128.000 163.000 ;
        RECT 109.000 157.000 115.000 158.000 ;
        RECT 118.000 158.000 121.000 162.000 ;
        RECT 125.000 161.000 127.000 162.000 ;
        RECT 125.000 160.000 126.000 161.000 ;
        RECT 118.000 157.000 129.000 158.000 ;
        RECT 110.000 156.000 117.000 157.000 ;
        RECT 118.000 156.000 130.000 157.000 ;
        RECT 110.000 155.000 116.000 156.000 ;
        RECT 109.000 154.000 115.000 155.000 ;
        RECT 109.000 153.000 111.000 154.000 ;
        RECT 108.000 152.000 111.000 153.000 ;
        RECT 107.000 151.000 111.000 152.000 ;
        RECT 106.000 150.000 110.000 151.000 ;
        RECT 112.000 150.000 115.000 154.000 ;
        RECT 120.000 153.000 121.000 154.000 ;
        RECT 119.000 152.000 121.000 153.000 ;
        RECT 118.000 150.000 121.000 152.000 ;
        RECT 125.000 150.000 128.000 156.000 ;
        RECT 106.000 149.000 109.000 150.000 ;
        RECT 112.000 149.000 114.000 150.000 ;
        RECT 118.000 149.000 127.000 150.000 ;
        RECT 107.000 148.000 108.000 149.000 ;
        RECT 112.000 148.000 113.000 149.000 ;
        RECT 118.000 148.000 126.000 149.000 ;
        RECT 68.100 137.300 89.700 140.000 ;
        RECT 68.100 134.600 92.400 137.300 ;
        RECT 62.700 129.200 97.800 134.600 ;
        RECT 60.000 118.400 100.500 129.200 ;
        RECT 60.000 115.700 68.100 118.400 ;
        RECT 60.000 113.000 65.400 115.700 ;
        RECT 62.700 110.300 65.400 113.000 ;
        RECT 76.200 110.300 84.300 118.400 ;
        RECT 92.400 115.700 100.500 118.400 ;
        RECT 95.100 113.000 100.500 115.700 ;
        RECT 95.100 110.300 97.800 113.000 ;
        RECT 62.700 107.600 68.100 110.300 ;
        RECT 73.500 107.600 87.000 110.300 ;
        RECT 92.400 107.600 97.800 110.300 ;
        RECT 65.400 104.900 78.900 107.600 ;
        RECT 81.600 104.900 97.800 107.600 ;
        RECT 65.400 102.200 76.200 104.900 ;
        RECT 84.300 102.200 92.400 104.900 ;
        RECT 70.800 96.800 89.700 102.200 ;
        RECT 54.600 94.100 57.300 96.800 ;
        RECT 70.800 94.100 73.500 96.800 ;
        RECT 76.200 94.100 78.900 96.800 ;
        RECT 81.600 94.100 84.300 96.800 ;
        RECT 87.000 94.100 89.700 96.800 ;
        RECT 103.200 94.100 105.900 96.800 ;
        RECT 51.900 91.400 60.000 94.100 ;
        RECT 100.500 91.400 108.600 94.100 ;
        RECT 51.900 88.700 62.700 91.400 ;
        RECT 97.800 88.700 108.600 91.400 ;
        RECT 51.900 86.000 68.100 88.700 ;
        RECT 92.400 86.000 108.600 88.700 ;
        RECT 51.900 83.300 73.500 86.000 ;
        RECT 87.000 83.300 105.900 86.000 ;
        RECT 68.100 80.600 78.900 83.300 ;
        RECT 81.600 80.600 92.400 83.300 ;
        RECT 73.500 75.200 87.000 80.600 ;
        RECT 68.100 72.500 78.900 75.200 ;
        RECT 81.600 72.500 92.400 75.200 ;
        RECT 62.700 69.800 73.500 72.500 ;
        RECT 87.000 69.800 97.800 72.500 ;
        RECT 54.600 67.100 70.800 69.800 ;
        RECT 89.700 67.100 105.900 69.800 ;
        RECT 51.900 61.700 65.400 67.100 ;
        RECT 95.100 61.700 108.600 67.100 ;
        RECT 54.600 59.000 62.700 61.700 ;
        RECT 70.800 59.000 73.500 61.700 ;
        RECT 76.200 59.000 78.900 61.700 ;
        RECT 81.600 59.000 84.300 61.700 ;
        RECT 87.000 59.000 89.700 61.700 ;
        RECT 97.800 59.000 105.900 61.700 ;
        RECT 70.800 53.600 89.700 59.000 ;
        RECT 65.400 50.900 76.200 53.600 ;
        RECT 84.300 50.900 92.400 53.600 ;
        RECT 65.400 48.200 78.900 50.900 ;
        RECT 81.600 48.200 97.800 50.900 ;
        RECT 62.700 45.500 68.100 48.200 ;
        RECT 73.500 45.500 87.000 48.200 ;
        RECT 92.400 45.500 97.800 48.200 ;
        RECT 62.700 42.800 65.400 45.500 ;
        RECT 60.000 40.100 65.400 42.800 ;
        RECT 60.000 37.400 68.100 40.100 ;
        RECT 76.200 37.400 84.300 45.500 ;
        RECT 95.100 42.800 97.800 45.500 ;
        RECT 95.100 40.100 100.500 42.800 ;
        RECT 92.400 37.400 100.500 40.100 ;
        RECT 60.000 26.600 100.500 37.400 ;
        RECT 62.700 21.200 97.800 26.600 ;
        RECT 68.100 18.500 92.400 21.200 ;
        RECT 68.100 15.800 89.700 18.500 ;
      LAYER met2 ;
        RECT 50.000 40.000 110.000 170.000 ;
        RECT 25.000 10.000 130.000 40.000 ;
      LAYER met3 ;
        RECT 50.000 40.000 110.000 170.000 ;
        RECT 25.000 10.000 130.000 40.000 ;
      LAYER met4 ;
        RECT 83.000 164.000 84.000 165.000 ;
        RECT 93.000 164.000 94.000 165.000 ;
        RECT 114.000 164.000 115.000 165.000 ;
        RECT 40.000 163.000 45.000 164.000 ;
        RECT 39.000 162.000 44.000 163.000 ;
        RECT 37.000 154.000 38.000 155.000 ;
        RECT 37.000 153.000 39.000 154.000 ;
        RECT 41.000 153.000 44.000 162.000 ;
        RECT 49.000 162.000 59.000 164.000 ;
        RECT 49.000 160.000 52.000 162.000 ;
        RECT 50.000 159.000 52.000 160.000 ;
        RECT 51.000 158.000 52.000 159.000 ;
        RECT 56.000 157.000 59.000 162.000 ;
        RECT 69.000 157.000 72.000 164.000 ;
        RECT 75.000 163.000 84.000 164.000 ;
        RECT 75.000 162.000 77.000 163.000 ;
        RECT 79.000 162.000 84.000 163.000 ;
        RECT 75.000 161.000 76.000 162.000 ;
        RECT 53.000 156.000 61.000 157.000 ;
        RECT 66.000 156.000 74.000 157.000 ;
        RECT 53.000 155.000 60.000 156.000 ;
        RECT 66.000 155.000 73.000 156.000 ;
        RECT 51.000 153.000 52.000 154.000 ;
        RECT 37.000 152.000 45.000 153.000 ;
        RECT 50.000 152.000 52.000 153.000 ;
        RECT 37.000 151.000 47.000 152.000 ;
        RECT 38.000 150.000 48.000 151.000 ;
        RECT 49.000 150.000 52.000 152.000 ;
        RECT 56.000 150.000 59.000 155.000 ;
        RECT 64.000 153.000 65.000 154.000 ;
        RECT 63.000 152.000 65.000 153.000 ;
        RECT 62.000 150.000 65.000 152.000 ;
        RECT 69.000 150.000 72.000 155.000 ;
        RECT 81.000 150.000 84.000 162.000 ;
        RECT 85.000 163.000 94.000 164.000 ;
        RECT 97.000 163.000 105.000 164.000 ;
        RECT 107.000 163.000 108.000 164.000 ;
        RECT 85.000 162.000 87.000 163.000 ;
        RECT 89.000 162.000 94.000 163.000 ;
        RECT 96.000 162.000 105.000 163.000 ;
        RECT 85.000 161.000 86.000 162.000 ;
        RECT 91.000 150.000 94.000 162.000 ;
        RECT 95.000 150.000 98.000 162.000 ;
        RECT 41.000 148.000 44.000 150.000 ;
        RECT 49.000 149.000 58.000 150.000 ;
        RECT 62.000 149.000 71.000 150.000 ;
        RECT 81.000 149.000 83.000 150.000 ;
        RECT 91.000 149.000 93.000 150.000 ;
        RECT 96.000 149.000 98.000 150.000 ;
        RECT 49.000 148.000 57.000 149.000 ;
        RECT 62.000 148.000 70.000 149.000 ;
        RECT 81.000 148.000 82.000 149.000 ;
        RECT 91.000 148.000 92.000 149.000 ;
        RECT 97.000 148.000 98.000 149.000 ;
        RECT 102.000 148.000 105.000 162.000 ;
        RECT 106.000 162.000 109.000 163.000 ;
        RECT 106.000 161.000 110.000 162.000 ;
        RECT 107.000 160.000 111.000 161.000 ;
        RECT 108.000 159.000 111.000 160.000 ;
        RECT 109.000 158.000 111.000 159.000 ;
        RECT 112.000 158.000 115.000 164.000 ;
        RECT 120.000 163.000 129.000 164.000 ;
        RECT 119.000 162.000 128.000 163.000 ;
        RECT 109.000 157.000 115.000 158.000 ;
        RECT 118.000 158.000 121.000 162.000 ;
        RECT 125.000 161.000 127.000 162.000 ;
        RECT 125.000 160.000 126.000 161.000 ;
        RECT 118.000 157.000 129.000 158.000 ;
        RECT 110.000 156.000 117.000 157.000 ;
        RECT 118.000 156.000 130.000 157.000 ;
        RECT 110.000 155.000 116.000 156.000 ;
        RECT 109.000 154.000 115.000 155.000 ;
        RECT 109.000 153.000 111.000 154.000 ;
        RECT 108.000 152.000 111.000 153.000 ;
        RECT 107.000 151.000 111.000 152.000 ;
        RECT 106.000 150.000 110.000 151.000 ;
        RECT 112.000 150.000 115.000 154.000 ;
        RECT 120.000 153.000 121.000 154.000 ;
        RECT 119.000 152.000 121.000 153.000 ;
        RECT 118.000 150.000 121.000 152.000 ;
        RECT 125.000 150.000 128.000 156.000 ;
        RECT 106.000 149.000 109.000 150.000 ;
        RECT 112.000 149.000 114.000 150.000 ;
        RECT 118.000 149.000 127.000 150.000 ;
        RECT 107.000 148.000 108.000 149.000 ;
        RECT 112.000 148.000 113.000 149.000 ;
        RECT 118.000 148.000 126.000 149.000 ;
        RECT 68.100 137.300 89.700 140.000 ;
        RECT 68.100 134.600 92.400 137.300 ;
        RECT 62.700 129.200 97.800 134.600 ;
        RECT 60.000 118.400 100.500 129.200 ;
        RECT 60.000 115.700 68.100 118.400 ;
        RECT 60.000 113.000 65.400 115.700 ;
        RECT 62.700 110.300 65.400 113.000 ;
        RECT 76.200 110.300 84.300 118.400 ;
        RECT 92.400 115.700 100.500 118.400 ;
        RECT 95.100 113.000 100.500 115.700 ;
        RECT 95.100 110.300 97.800 113.000 ;
        RECT 62.700 107.600 68.100 110.300 ;
        RECT 73.500 107.600 87.000 110.300 ;
        RECT 92.400 107.600 97.800 110.300 ;
        RECT 65.400 104.900 78.900 107.600 ;
        RECT 81.600 104.900 97.800 107.600 ;
        RECT 65.400 102.200 76.200 104.900 ;
        RECT 84.300 102.200 92.400 104.900 ;
        RECT 70.800 96.800 89.700 102.200 ;
        RECT 54.600 94.100 57.300 96.800 ;
        RECT 70.800 94.100 73.500 96.800 ;
        RECT 76.200 94.100 78.900 96.800 ;
        RECT 81.600 94.100 84.300 96.800 ;
        RECT 87.000 94.100 89.700 96.800 ;
        RECT 103.200 94.100 105.900 96.800 ;
        RECT 51.900 91.400 60.000 94.100 ;
        RECT 100.500 91.400 108.600 94.100 ;
        RECT 51.900 88.700 62.700 91.400 ;
        RECT 97.800 88.700 108.600 91.400 ;
        RECT 51.900 86.000 68.100 88.700 ;
        RECT 92.400 86.000 108.600 88.700 ;
        RECT 51.900 83.300 73.500 86.000 ;
        RECT 87.000 83.300 105.900 86.000 ;
        RECT 68.100 80.600 78.900 83.300 ;
        RECT 81.600 80.600 92.400 83.300 ;
        RECT 73.500 75.200 87.000 80.600 ;
        RECT 68.100 72.500 78.900 75.200 ;
        RECT 81.600 72.500 92.400 75.200 ;
        RECT 62.700 69.800 73.500 72.500 ;
        RECT 87.000 69.800 97.800 72.500 ;
        RECT 54.600 67.100 70.800 69.800 ;
        RECT 89.700 67.100 105.900 69.800 ;
        RECT 51.900 61.700 65.400 67.100 ;
        RECT 95.100 61.700 108.600 67.100 ;
        RECT 54.600 59.000 62.700 61.700 ;
        RECT 70.800 59.000 73.500 61.700 ;
        RECT 76.200 59.000 78.900 61.700 ;
        RECT 81.600 59.000 84.300 61.700 ;
        RECT 87.000 59.000 89.700 61.700 ;
        RECT 97.800 59.000 105.900 61.700 ;
        RECT 70.800 53.600 89.700 59.000 ;
        RECT 65.400 50.900 76.200 53.600 ;
        RECT 84.300 50.900 92.400 53.600 ;
        RECT 65.400 48.200 78.900 50.900 ;
        RECT 81.600 48.200 97.800 50.900 ;
        RECT 62.700 45.500 68.100 48.200 ;
        RECT 73.500 45.500 87.000 48.200 ;
        RECT 92.400 45.500 97.800 48.200 ;
        RECT 62.700 42.800 65.400 45.500 ;
        RECT 60.000 40.100 65.400 42.800 ;
        RECT 60.000 37.400 68.100 40.100 ;
        RECT 76.200 37.400 84.300 45.500 ;
        RECT 95.100 42.800 97.800 45.500 ;
        RECT 95.100 40.100 100.500 42.800 ;
        RECT 92.400 37.400 100.500 40.100 ;
        RECT 60.000 26.600 100.500 37.400 ;
        RECT 62.700 21.200 97.800 26.600 ;
        RECT 68.100 18.500 92.400 21.200 ;
        RECT 68.100 15.800 89.700 18.500 ;
  END
END skullart
END LIBRARY

