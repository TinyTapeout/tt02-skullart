module user_project_wrapper (user_clock2,
    vccd1,
    vccd2,
    vdda1,
    vdda2,
    vssa1,
    vssa2,
    vssd1,
    vssd2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input vccd1;
 input vccd2;
 input vdda1;
 input vdda2;
 input vssa1;
 input vssa2;
 input vssd1;
 input vssd2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire sc_clk_in;
 wire sc_clk_out;
 wire sc_data_in;
 wire sc_data_out;
 wire sc_latch_out;
 wire sc_scan_out;
 wire sw_000_clk_out;
 wire sw_000_data_out;
 wire sw_000_latch_out;
 wire \sw_000_module_data_in[0] ;
 wire \sw_000_module_data_in[1] ;
 wire \sw_000_module_data_in[2] ;
 wire \sw_000_module_data_in[3] ;
 wire \sw_000_module_data_in[4] ;
 wire \sw_000_module_data_in[5] ;
 wire \sw_000_module_data_in[6] ;
 wire \sw_000_module_data_in[7] ;
 wire \sw_000_module_data_out[0] ;
 wire \sw_000_module_data_out[1] ;
 wire \sw_000_module_data_out[2] ;
 wire \sw_000_module_data_out[3] ;
 wire \sw_000_module_data_out[4] ;
 wire \sw_000_module_data_out[5] ;
 wire \sw_000_module_data_out[6] ;
 wire \sw_000_module_data_out[7] ;
 wire sw_000_scan_out;
 wire sw_001_clk_out;
 wire sw_001_data_out;
 wire sw_001_latch_out;
 wire \sw_001_module_data_in[0] ;
 wire \sw_001_module_data_in[1] ;
 wire \sw_001_module_data_in[2] ;
 wire \sw_001_module_data_in[3] ;
 wire \sw_001_module_data_in[4] ;
 wire \sw_001_module_data_in[5] ;
 wire \sw_001_module_data_in[6] ;
 wire \sw_001_module_data_in[7] ;
 wire \sw_001_module_data_out[0] ;
 wire \sw_001_module_data_out[1] ;
 wire \sw_001_module_data_out[2] ;
 wire \sw_001_module_data_out[3] ;
 wire \sw_001_module_data_out[4] ;
 wire \sw_001_module_data_out[5] ;
 wire \sw_001_module_data_out[6] ;
 wire \sw_001_module_data_out[7] ;
 wire sw_001_scan_out;
 wire sw_002_clk_out;
 wire sw_002_data_out;
 wire sw_002_latch_out;
 wire \sw_002_module_data_in[0] ;
 wire \sw_002_module_data_in[1] ;
 wire \sw_002_module_data_in[2] ;
 wire \sw_002_module_data_in[3] ;
 wire \sw_002_module_data_in[4] ;
 wire \sw_002_module_data_in[5] ;
 wire \sw_002_module_data_in[6] ;
 wire \sw_002_module_data_in[7] ;
 wire \sw_002_module_data_out[0] ;
 wire \sw_002_module_data_out[1] ;
 wire \sw_002_module_data_out[2] ;
 wire \sw_002_module_data_out[3] ;
 wire \sw_002_module_data_out[4] ;
 wire \sw_002_module_data_out[5] ;
 wire \sw_002_module_data_out[6] ;
 wire \sw_002_module_data_out[7] ;
 wire sw_002_scan_out;
 wire sw_003_clk_out;
 wire sw_003_data_out;
 wire sw_003_latch_out;
 wire \sw_003_module_data_in[0] ;
 wire \sw_003_module_data_in[1] ;
 wire \sw_003_module_data_in[2] ;
 wire \sw_003_module_data_in[3] ;
 wire \sw_003_module_data_in[4] ;
 wire \sw_003_module_data_in[5] ;
 wire \sw_003_module_data_in[6] ;
 wire \sw_003_module_data_in[7] ;
 wire \sw_003_module_data_out[0] ;
 wire \sw_003_module_data_out[1] ;
 wire \sw_003_module_data_out[2] ;
 wire \sw_003_module_data_out[3] ;
 wire \sw_003_module_data_out[4] ;
 wire \sw_003_module_data_out[5] ;
 wire \sw_003_module_data_out[6] ;
 wire \sw_003_module_data_out[7] ;
 wire sw_003_scan_out;
 wire sw_004_clk_out;
 wire sw_004_data_out;
 wire sw_004_latch_out;
 wire \sw_004_module_data_in[0] ;
 wire \sw_004_module_data_in[1] ;
 wire \sw_004_module_data_in[2] ;
 wire \sw_004_module_data_in[3] ;
 wire \sw_004_module_data_in[4] ;
 wire \sw_004_module_data_in[5] ;
 wire \sw_004_module_data_in[6] ;
 wire \sw_004_module_data_in[7] ;
 wire \sw_004_module_data_out[0] ;
 wire \sw_004_module_data_out[1] ;
 wire \sw_004_module_data_out[2] ;
 wire \sw_004_module_data_out[3] ;
 wire \sw_004_module_data_out[4] ;
 wire \sw_004_module_data_out[5] ;
 wire \sw_004_module_data_out[6] ;
 wire \sw_004_module_data_out[7] ;
 wire sw_004_scan_out;
 wire sw_005_clk_out;
 wire sw_005_data_out;
 wire sw_005_latch_out;
 wire \sw_005_module_data_in[0] ;
 wire \sw_005_module_data_in[1] ;
 wire \sw_005_module_data_in[2] ;
 wire \sw_005_module_data_in[3] ;
 wire \sw_005_module_data_in[4] ;
 wire \sw_005_module_data_in[5] ;
 wire \sw_005_module_data_in[6] ;
 wire \sw_005_module_data_in[7] ;
 wire \sw_005_module_data_out[0] ;
 wire \sw_005_module_data_out[1] ;
 wire \sw_005_module_data_out[2] ;
 wire \sw_005_module_data_out[3] ;
 wire \sw_005_module_data_out[4] ;
 wire \sw_005_module_data_out[5] ;
 wire \sw_005_module_data_out[6] ;
 wire \sw_005_module_data_out[7] ;
 wire sw_005_scan_out;
 wire sw_006_clk_out;
 wire sw_006_data_out;
 wire sw_006_latch_out;
 wire \sw_006_module_data_in[0] ;
 wire \sw_006_module_data_in[1] ;
 wire \sw_006_module_data_in[2] ;
 wire \sw_006_module_data_in[3] ;
 wire \sw_006_module_data_in[4] ;
 wire \sw_006_module_data_in[5] ;
 wire \sw_006_module_data_in[6] ;
 wire \sw_006_module_data_in[7] ;
 wire \sw_006_module_data_out[0] ;
 wire \sw_006_module_data_out[1] ;
 wire \sw_006_module_data_out[2] ;
 wire \sw_006_module_data_out[3] ;
 wire \sw_006_module_data_out[4] ;
 wire \sw_006_module_data_out[5] ;
 wire \sw_006_module_data_out[6] ;
 wire \sw_006_module_data_out[7] ;
 wire sw_006_scan_out;
 wire sw_007_clk_out;
 wire sw_007_data_out;
 wire sw_007_latch_out;
 wire \sw_007_module_data_in[0] ;
 wire \sw_007_module_data_in[1] ;
 wire \sw_007_module_data_in[2] ;
 wire \sw_007_module_data_in[3] ;
 wire \sw_007_module_data_in[4] ;
 wire \sw_007_module_data_in[5] ;
 wire \sw_007_module_data_in[6] ;
 wire \sw_007_module_data_in[7] ;
 wire \sw_007_module_data_out[0] ;
 wire \sw_007_module_data_out[1] ;
 wire \sw_007_module_data_out[2] ;
 wire \sw_007_module_data_out[3] ;
 wire \sw_007_module_data_out[4] ;
 wire \sw_007_module_data_out[5] ;
 wire \sw_007_module_data_out[6] ;
 wire \sw_007_module_data_out[7] ;
 wire sw_007_scan_out;
 wire sw_008_clk_out;
 wire sw_008_data_out;
 wire sw_008_latch_out;
 wire \sw_008_module_data_in[0] ;
 wire \sw_008_module_data_in[1] ;
 wire \sw_008_module_data_in[2] ;
 wire \sw_008_module_data_in[3] ;
 wire \sw_008_module_data_in[4] ;
 wire \sw_008_module_data_in[5] ;
 wire \sw_008_module_data_in[6] ;
 wire \sw_008_module_data_in[7] ;
 wire \sw_008_module_data_out[0] ;
 wire \sw_008_module_data_out[1] ;
 wire \sw_008_module_data_out[2] ;
 wire \sw_008_module_data_out[3] ;
 wire \sw_008_module_data_out[4] ;
 wire \sw_008_module_data_out[5] ;
 wire \sw_008_module_data_out[6] ;
 wire \sw_008_module_data_out[7] ;
 wire sw_008_scan_out;
 wire sw_009_clk_out;
 wire sw_009_data_out;
 wire sw_009_latch_out;
 wire \sw_009_module_data_in[0] ;
 wire \sw_009_module_data_in[1] ;
 wire \sw_009_module_data_in[2] ;
 wire \sw_009_module_data_in[3] ;
 wire \sw_009_module_data_in[4] ;
 wire \sw_009_module_data_in[5] ;
 wire \sw_009_module_data_in[6] ;
 wire \sw_009_module_data_in[7] ;
 wire \sw_009_module_data_out[0] ;
 wire \sw_009_module_data_out[1] ;
 wire \sw_009_module_data_out[2] ;
 wire \sw_009_module_data_out[3] ;
 wire \sw_009_module_data_out[4] ;
 wire \sw_009_module_data_out[5] ;
 wire \sw_009_module_data_out[6] ;
 wire \sw_009_module_data_out[7] ;
 wire sw_009_scan_out;
 wire sw_010_clk_out;
 wire sw_010_data_out;
 wire sw_010_latch_out;
 wire \sw_010_module_data_in[0] ;
 wire \sw_010_module_data_in[1] ;
 wire \sw_010_module_data_in[2] ;
 wire \sw_010_module_data_in[3] ;
 wire \sw_010_module_data_in[4] ;
 wire \sw_010_module_data_in[5] ;
 wire \sw_010_module_data_in[6] ;
 wire \sw_010_module_data_in[7] ;
 wire \sw_010_module_data_out[0] ;
 wire \sw_010_module_data_out[1] ;
 wire \sw_010_module_data_out[2] ;
 wire \sw_010_module_data_out[3] ;
 wire \sw_010_module_data_out[4] ;
 wire \sw_010_module_data_out[5] ;
 wire \sw_010_module_data_out[6] ;
 wire \sw_010_module_data_out[7] ;
 wire sw_010_scan_out;
 wire sw_011_clk_out;
 wire sw_011_data_out;
 wire sw_011_latch_out;
 wire \sw_011_module_data_in[0] ;
 wire \sw_011_module_data_in[1] ;
 wire \sw_011_module_data_in[2] ;
 wire \sw_011_module_data_in[3] ;
 wire \sw_011_module_data_in[4] ;
 wire \sw_011_module_data_in[5] ;
 wire \sw_011_module_data_in[6] ;
 wire \sw_011_module_data_in[7] ;
 wire \sw_011_module_data_out[0] ;
 wire \sw_011_module_data_out[1] ;
 wire \sw_011_module_data_out[2] ;
 wire \sw_011_module_data_out[3] ;
 wire \sw_011_module_data_out[4] ;
 wire \sw_011_module_data_out[5] ;
 wire \sw_011_module_data_out[6] ;
 wire \sw_011_module_data_out[7] ;
 wire sw_011_scan_out;
 wire sw_012_clk_out;
 wire sw_012_data_out;
 wire sw_012_latch_out;
 wire \sw_012_module_data_in[0] ;
 wire \sw_012_module_data_in[1] ;
 wire \sw_012_module_data_in[2] ;
 wire \sw_012_module_data_in[3] ;
 wire \sw_012_module_data_in[4] ;
 wire \sw_012_module_data_in[5] ;
 wire \sw_012_module_data_in[6] ;
 wire \sw_012_module_data_in[7] ;
 wire \sw_012_module_data_out[0] ;
 wire \sw_012_module_data_out[1] ;
 wire \sw_012_module_data_out[2] ;
 wire \sw_012_module_data_out[3] ;
 wire \sw_012_module_data_out[4] ;
 wire \sw_012_module_data_out[5] ;
 wire \sw_012_module_data_out[6] ;
 wire \sw_012_module_data_out[7] ;
 wire sw_012_scan_out;
 wire sw_013_clk_out;
 wire sw_013_data_out;
 wire sw_013_latch_out;
 wire \sw_013_module_data_in[0] ;
 wire \sw_013_module_data_in[1] ;
 wire \sw_013_module_data_in[2] ;
 wire \sw_013_module_data_in[3] ;
 wire \sw_013_module_data_in[4] ;
 wire \sw_013_module_data_in[5] ;
 wire \sw_013_module_data_in[6] ;
 wire \sw_013_module_data_in[7] ;
 wire \sw_013_module_data_out[0] ;
 wire \sw_013_module_data_out[1] ;
 wire \sw_013_module_data_out[2] ;
 wire \sw_013_module_data_out[3] ;
 wire \sw_013_module_data_out[4] ;
 wire \sw_013_module_data_out[5] ;
 wire \sw_013_module_data_out[6] ;
 wire \sw_013_module_data_out[7] ;
 wire sw_013_scan_out;
 wire sw_014_clk_out;
 wire sw_014_data_out;
 wire sw_014_latch_out;
 wire \sw_014_module_data_in[0] ;
 wire \sw_014_module_data_in[1] ;
 wire \sw_014_module_data_in[2] ;
 wire \sw_014_module_data_in[3] ;
 wire \sw_014_module_data_in[4] ;
 wire \sw_014_module_data_in[5] ;
 wire \sw_014_module_data_in[6] ;
 wire \sw_014_module_data_in[7] ;
 wire \sw_014_module_data_out[0] ;
 wire \sw_014_module_data_out[1] ;
 wire \sw_014_module_data_out[2] ;
 wire \sw_014_module_data_out[3] ;
 wire \sw_014_module_data_out[4] ;
 wire \sw_014_module_data_out[5] ;
 wire \sw_014_module_data_out[6] ;
 wire \sw_014_module_data_out[7] ;
 wire sw_014_scan_out;
 wire sw_015_clk_out;
 wire sw_015_data_out;
 wire sw_015_latch_out;
 wire \sw_015_module_data_in[0] ;
 wire \sw_015_module_data_in[1] ;
 wire \sw_015_module_data_in[2] ;
 wire \sw_015_module_data_in[3] ;
 wire \sw_015_module_data_in[4] ;
 wire \sw_015_module_data_in[5] ;
 wire \sw_015_module_data_in[6] ;
 wire \sw_015_module_data_in[7] ;
 wire \sw_015_module_data_out[0] ;
 wire \sw_015_module_data_out[1] ;
 wire \sw_015_module_data_out[2] ;
 wire \sw_015_module_data_out[3] ;
 wire \sw_015_module_data_out[4] ;
 wire \sw_015_module_data_out[5] ;
 wire \sw_015_module_data_out[6] ;
 wire \sw_015_module_data_out[7] ;
 wire sw_015_scan_out;
 wire sw_016_clk_out;
 wire sw_016_data_out;
 wire sw_016_latch_out;
 wire \sw_016_module_data_in[0] ;
 wire \sw_016_module_data_in[1] ;
 wire \sw_016_module_data_in[2] ;
 wire \sw_016_module_data_in[3] ;
 wire \sw_016_module_data_in[4] ;
 wire \sw_016_module_data_in[5] ;
 wire \sw_016_module_data_in[6] ;
 wire \sw_016_module_data_in[7] ;
 wire \sw_016_module_data_out[0] ;
 wire \sw_016_module_data_out[1] ;
 wire \sw_016_module_data_out[2] ;
 wire \sw_016_module_data_out[3] ;
 wire \sw_016_module_data_out[4] ;
 wire \sw_016_module_data_out[5] ;
 wire \sw_016_module_data_out[6] ;
 wire \sw_016_module_data_out[7] ;
 wire sw_016_scan_out;
 wire sw_017_clk_out;
 wire sw_017_data_out;
 wire sw_017_latch_out;
 wire \sw_017_module_data_in[0] ;
 wire \sw_017_module_data_in[1] ;
 wire \sw_017_module_data_in[2] ;
 wire \sw_017_module_data_in[3] ;
 wire \sw_017_module_data_in[4] ;
 wire \sw_017_module_data_in[5] ;
 wire \sw_017_module_data_in[6] ;
 wire \sw_017_module_data_in[7] ;
 wire \sw_017_module_data_out[0] ;
 wire \sw_017_module_data_out[1] ;
 wire \sw_017_module_data_out[2] ;
 wire \sw_017_module_data_out[3] ;
 wire \sw_017_module_data_out[4] ;
 wire \sw_017_module_data_out[5] ;
 wire \sw_017_module_data_out[6] ;
 wire \sw_017_module_data_out[7] ;
 wire sw_017_scan_out;
 wire sw_018_clk_out;
 wire sw_018_data_out;
 wire sw_018_latch_out;
 wire \sw_018_module_data_in[0] ;
 wire \sw_018_module_data_in[1] ;
 wire \sw_018_module_data_in[2] ;
 wire \sw_018_module_data_in[3] ;
 wire \sw_018_module_data_in[4] ;
 wire \sw_018_module_data_in[5] ;
 wire \sw_018_module_data_in[6] ;
 wire \sw_018_module_data_in[7] ;
 wire \sw_018_module_data_out[0] ;
 wire \sw_018_module_data_out[1] ;
 wire \sw_018_module_data_out[2] ;
 wire \sw_018_module_data_out[3] ;
 wire \sw_018_module_data_out[4] ;
 wire \sw_018_module_data_out[5] ;
 wire \sw_018_module_data_out[6] ;
 wire \sw_018_module_data_out[7] ;
 wire sw_018_scan_out;
 wire sw_019_clk_out;
 wire sw_019_data_out;
 wire sw_019_latch_out;
 wire \sw_019_module_data_in[0] ;
 wire \sw_019_module_data_in[1] ;
 wire \sw_019_module_data_in[2] ;
 wire \sw_019_module_data_in[3] ;
 wire \sw_019_module_data_in[4] ;
 wire \sw_019_module_data_in[5] ;
 wire \sw_019_module_data_in[6] ;
 wire \sw_019_module_data_in[7] ;
 wire \sw_019_module_data_out[0] ;
 wire \sw_019_module_data_out[1] ;
 wire \sw_019_module_data_out[2] ;
 wire \sw_019_module_data_out[3] ;
 wire \sw_019_module_data_out[4] ;
 wire \sw_019_module_data_out[5] ;
 wire \sw_019_module_data_out[6] ;
 wire \sw_019_module_data_out[7] ;
 wire sw_019_scan_out;
 wire sw_020_clk_out;
 wire sw_020_data_out;
 wire sw_020_latch_out;
 wire \sw_020_module_data_in[0] ;
 wire \sw_020_module_data_in[1] ;
 wire \sw_020_module_data_in[2] ;
 wire \sw_020_module_data_in[3] ;
 wire \sw_020_module_data_in[4] ;
 wire \sw_020_module_data_in[5] ;
 wire \sw_020_module_data_in[6] ;
 wire \sw_020_module_data_in[7] ;
 wire \sw_020_module_data_out[0] ;
 wire \sw_020_module_data_out[1] ;
 wire \sw_020_module_data_out[2] ;
 wire \sw_020_module_data_out[3] ;
 wire \sw_020_module_data_out[4] ;
 wire \sw_020_module_data_out[5] ;
 wire \sw_020_module_data_out[6] ;
 wire \sw_020_module_data_out[7] ;
 wire sw_020_scan_out;
 wire sw_021_clk_out;
 wire sw_021_data_out;
 wire sw_021_latch_out;
 wire \sw_021_module_data_in[0] ;
 wire \sw_021_module_data_in[1] ;
 wire \sw_021_module_data_in[2] ;
 wire \sw_021_module_data_in[3] ;
 wire \sw_021_module_data_in[4] ;
 wire \sw_021_module_data_in[5] ;
 wire \sw_021_module_data_in[6] ;
 wire \sw_021_module_data_in[7] ;
 wire \sw_021_module_data_out[0] ;
 wire \sw_021_module_data_out[1] ;
 wire \sw_021_module_data_out[2] ;
 wire \sw_021_module_data_out[3] ;
 wire \sw_021_module_data_out[4] ;
 wire \sw_021_module_data_out[5] ;
 wire \sw_021_module_data_out[6] ;
 wire \sw_021_module_data_out[7] ;
 wire sw_021_scan_out;
 wire sw_022_clk_out;
 wire sw_022_data_out;
 wire sw_022_latch_out;
 wire \sw_022_module_data_in[0] ;
 wire \sw_022_module_data_in[1] ;
 wire \sw_022_module_data_in[2] ;
 wire \sw_022_module_data_in[3] ;
 wire \sw_022_module_data_in[4] ;
 wire \sw_022_module_data_in[5] ;
 wire \sw_022_module_data_in[6] ;
 wire \sw_022_module_data_in[7] ;
 wire \sw_022_module_data_out[0] ;
 wire \sw_022_module_data_out[1] ;
 wire \sw_022_module_data_out[2] ;
 wire \sw_022_module_data_out[3] ;
 wire \sw_022_module_data_out[4] ;
 wire \sw_022_module_data_out[5] ;
 wire \sw_022_module_data_out[6] ;
 wire \sw_022_module_data_out[7] ;
 wire sw_022_scan_out;
 wire sw_023_clk_out;
 wire sw_023_data_out;
 wire sw_023_latch_out;
 wire \sw_023_module_data_in[0] ;
 wire \sw_023_module_data_in[1] ;
 wire \sw_023_module_data_in[2] ;
 wire \sw_023_module_data_in[3] ;
 wire \sw_023_module_data_in[4] ;
 wire \sw_023_module_data_in[5] ;
 wire \sw_023_module_data_in[6] ;
 wire \sw_023_module_data_in[7] ;
 wire \sw_023_module_data_out[0] ;
 wire \sw_023_module_data_out[1] ;
 wire \sw_023_module_data_out[2] ;
 wire \sw_023_module_data_out[3] ;
 wire \sw_023_module_data_out[4] ;
 wire \sw_023_module_data_out[5] ;
 wire \sw_023_module_data_out[6] ;
 wire \sw_023_module_data_out[7] ;
 wire sw_023_scan_out;
 wire sw_024_clk_out;
 wire sw_024_data_out;
 wire sw_024_latch_out;
 wire \sw_024_module_data_in[0] ;
 wire \sw_024_module_data_in[1] ;
 wire \sw_024_module_data_in[2] ;
 wire \sw_024_module_data_in[3] ;
 wire \sw_024_module_data_in[4] ;
 wire \sw_024_module_data_in[5] ;
 wire \sw_024_module_data_in[6] ;
 wire \sw_024_module_data_in[7] ;
 wire \sw_024_module_data_out[0] ;
 wire \sw_024_module_data_out[1] ;
 wire \sw_024_module_data_out[2] ;
 wire \sw_024_module_data_out[3] ;
 wire \sw_024_module_data_out[4] ;
 wire \sw_024_module_data_out[5] ;
 wire \sw_024_module_data_out[6] ;
 wire \sw_024_module_data_out[7] ;
 wire sw_024_scan_out;
 wire sw_025_clk_out;
 wire sw_025_data_out;
 wire sw_025_latch_out;
 wire \sw_025_module_data_in[0] ;
 wire \sw_025_module_data_in[1] ;
 wire \sw_025_module_data_in[2] ;
 wire \sw_025_module_data_in[3] ;
 wire \sw_025_module_data_in[4] ;
 wire \sw_025_module_data_in[5] ;
 wire \sw_025_module_data_in[6] ;
 wire \sw_025_module_data_in[7] ;
 wire \sw_025_module_data_out[0] ;
 wire \sw_025_module_data_out[1] ;
 wire \sw_025_module_data_out[2] ;
 wire \sw_025_module_data_out[3] ;
 wire \sw_025_module_data_out[4] ;
 wire \sw_025_module_data_out[5] ;
 wire \sw_025_module_data_out[6] ;
 wire \sw_025_module_data_out[7] ;
 wire sw_025_scan_out;
 wire sw_026_clk_out;
 wire sw_026_data_out;
 wire sw_026_latch_out;
 wire \sw_026_module_data_in[0] ;
 wire \sw_026_module_data_in[1] ;
 wire \sw_026_module_data_in[2] ;
 wire \sw_026_module_data_in[3] ;
 wire \sw_026_module_data_in[4] ;
 wire \sw_026_module_data_in[5] ;
 wire \sw_026_module_data_in[6] ;
 wire \sw_026_module_data_in[7] ;
 wire \sw_026_module_data_out[0] ;
 wire \sw_026_module_data_out[1] ;
 wire \sw_026_module_data_out[2] ;
 wire \sw_026_module_data_out[3] ;
 wire \sw_026_module_data_out[4] ;
 wire \sw_026_module_data_out[5] ;
 wire \sw_026_module_data_out[6] ;
 wire \sw_026_module_data_out[7] ;
 wire sw_026_scan_out;
 wire sw_027_clk_out;
 wire sw_027_data_out;
 wire sw_027_latch_out;
 wire \sw_027_module_data_in[0] ;
 wire \sw_027_module_data_in[1] ;
 wire \sw_027_module_data_in[2] ;
 wire \sw_027_module_data_in[3] ;
 wire \sw_027_module_data_in[4] ;
 wire \sw_027_module_data_in[5] ;
 wire \sw_027_module_data_in[6] ;
 wire \sw_027_module_data_in[7] ;
 wire \sw_027_module_data_out[0] ;
 wire \sw_027_module_data_out[1] ;
 wire \sw_027_module_data_out[2] ;
 wire \sw_027_module_data_out[3] ;
 wire \sw_027_module_data_out[4] ;
 wire \sw_027_module_data_out[5] ;
 wire \sw_027_module_data_out[6] ;
 wire \sw_027_module_data_out[7] ;
 wire sw_027_scan_out;
 wire sw_028_clk_out;
 wire sw_028_data_out;
 wire sw_028_latch_out;
 wire \sw_028_module_data_in[0] ;
 wire \sw_028_module_data_in[1] ;
 wire \sw_028_module_data_in[2] ;
 wire \sw_028_module_data_in[3] ;
 wire \sw_028_module_data_in[4] ;
 wire \sw_028_module_data_in[5] ;
 wire \sw_028_module_data_in[6] ;
 wire \sw_028_module_data_in[7] ;
 wire \sw_028_module_data_out[0] ;
 wire \sw_028_module_data_out[1] ;
 wire \sw_028_module_data_out[2] ;
 wire \sw_028_module_data_out[3] ;
 wire \sw_028_module_data_out[4] ;
 wire \sw_028_module_data_out[5] ;
 wire \sw_028_module_data_out[6] ;
 wire \sw_028_module_data_out[7] ;
 wire sw_028_scan_out;
 wire sw_029_clk_out;
 wire sw_029_data_out;
 wire sw_029_latch_out;
 wire \sw_029_module_data_in[0] ;
 wire \sw_029_module_data_in[1] ;
 wire \sw_029_module_data_in[2] ;
 wire \sw_029_module_data_in[3] ;
 wire \sw_029_module_data_in[4] ;
 wire \sw_029_module_data_in[5] ;
 wire \sw_029_module_data_in[6] ;
 wire \sw_029_module_data_in[7] ;
 wire \sw_029_module_data_out[0] ;
 wire \sw_029_module_data_out[1] ;
 wire \sw_029_module_data_out[2] ;
 wire \sw_029_module_data_out[3] ;
 wire \sw_029_module_data_out[4] ;
 wire \sw_029_module_data_out[5] ;
 wire \sw_029_module_data_out[6] ;
 wire \sw_029_module_data_out[7] ;
 wire sw_029_scan_out;
 wire sw_030_clk_out;
 wire sw_030_data_out;
 wire sw_030_latch_out;
 wire \sw_030_module_data_in[0] ;
 wire \sw_030_module_data_in[1] ;
 wire \sw_030_module_data_in[2] ;
 wire \sw_030_module_data_in[3] ;
 wire \sw_030_module_data_in[4] ;
 wire \sw_030_module_data_in[5] ;
 wire \sw_030_module_data_in[6] ;
 wire \sw_030_module_data_in[7] ;
 wire \sw_030_module_data_out[0] ;
 wire \sw_030_module_data_out[1] ;
 wire \sw_030_module_data_out[2] ;
 wire \sw_030_module_data_out[3] ;
 wire \sw_030_module_data_out[4] ;
 wire \sw_030_module_data_out[5] ;
 wire \sw_030_module_data_out[6] ;
 wire \sw_030_module_data_out[7] ;
 wire sw_030_scan_out;
 wire sw_031_clk_out;
 wire sw_031_data_out;
 wire sw_031_latch_out;
 wire \sw_031_module_data_in[0] ;
 wire \sw_031_module_data_in[1] ;
 wire \sw_031_module_data_in[2] ;
 wire \sw_031_module_data_in[3] ;
 wire \sw_031_module_data_in[4] ;
 wire \sw_031_module_data_in[5] ;
 wire \sw_031_module_data_in[6] ;
 wire \sw_031_module_data_in[7] ;
 wire \sw_031_module_data_out[0] ;
 wire \sw_031_module_data_out[1] ;
 wire \sw_031_module_data_out[2] ;
 wire \sw_031_module_data_out[3] ;
 wire \sw_031_module_data_out[4] ;
 wire \sw_031_module_data_out[5] ;
 wire \sw_031_module_data_out[6] ;
 wire \sw_031_module_data_out[7] ;
 wire sw_031_scan_out;
 wire sw_032_clk_out;
 wire sw_032_data_out;
 wire sw_032_latch_out;
 wire \sw_032_module_data_in[0] ;
 wire \sw_032_module_data_in[1] ;
 wire \sw_032_module_data_in[2] ;
 wire \sw_032_module_data_in[3] ;
 wire \sw_032_module_data_in[4] ;
 wire \sw_032_module_data_in[5] ;
 wire \sw_032_module_data_in[6] ;
 wire \sw_032_module_data_in[7] ;
 wire \sw_032_module_data_out[0] ;
 wire \sw_032_module_data_out[1] ;
 wire \sw_032_module_data_out[2] ;
 wire \sw_032_module_data_out[3] ;
 wire \sw_032_module_data_out[4] ;
 wire \sw_032_module_data_out[5] ;
 wire \sw_032_module_data_out[6] ;
 wire \sw_032_module_data_out[7] ;
 wire sw_032_scan_out;
 wire sw_033_clk_out;
 wire sw_033_data_out;
 wire sw_033_latch_out;
 wire \sw_033_module_data_in[0] ;
 wire \sw_033_module_data_in[1] ;
 wire \sw_033_module_data_in[2] ;
 wire \sw_033_module_data_in[3] ;
 wire \sw_033_module_data_in[4] ;
 wire \sw_033_module_data_in[5] ;
 wire \sw_033_module_data_in[6] ;
 wire \sw_033_module_data_in[7] ;
 wire \sw_033_module_data_out[0] ;
 wire \sw_033_module_data_out[1] ;
 wire \sw_033_module_data_out[2] ;
 wire \sw_033_module_data_out[3] ;
 wire \sw_033_module_data_out[4] ;
 wire \sw_033_module_data_out[5] ;
 wire \sw_033_module_data_out[6] ;
 wire \sw_033_module_data_out[7] ;
 wire sw_033_scan_out;
 wire sw_034_clk_out;
 wire sw_034_data_out;
 wire sw_034_latch_out;
 wire \sw_034_module_data_in[0] ;
 wire \sw_034_module_data_in[1] ;
 wire \sw_034_module_data_in[2] ;
 wire \sw_034_module_data_in[3] ;
 wire \sw_034_module_data_in[4] ;
 wire \sw_034_module_data_in[5] ;
 wire \sw_034_module_data_in[6] ;
 wire \sw_034_module_data_in[7] ;
 wire \sw_034_module_data_out[0] ;
 wire \sw_034_module_data_out[1] ;
 wire \sw_034_module_data_out[2] ;
 wire \sw_034_module_data_out[3] ;
 wire \sw_034_module_data_out[4] ;
 wire \sw_034_module_data_out[5] ;
 wire \sw_034_module_data_out[6] ;
 wire \sw_034_module_data_out[7] ;
 wire sw_034_scan_out;
 wire sw_035_clk_out;
 wire sw_035_data_out;
 wire sw_035_latch_out;
 wire \sw_035_module_data_in[0] ;
 wire \sw_035_module_data_in[1] ;
 wire \sw_035_module_data_in[2] ;
 wire \sw_035_module_data_in[3] ;
 wire \sw_035_module_data_in[4] ;
 wire \sw_035_module_data_in[5] ;
 wire \sw_035_module_data_in[6] ;
 wire \sw_035_module_data_in[7] ;
 wire \sw_035_module_data_out[0] ;
 wire \sw_035_module_data_out[1] ;
 wire \sw_035_module_data_out[2] ;
 wire \sw_035_module_data_out[3] ;
 wire \sw_035_module_data_out[4] ;
 wire \sw_035_module_data_out[5] ;
 wire \sw_035_module_data_out[6] ;
 wire \sw_035_module_data_out[7] ;
 wire sw_035_scan_out;
 wire sw_036_clk_out;
 wire sw_036_data_out;
 wire sw_036_latch_out;
 wire \sw_036_module_data_in[0] ;
 wire \sw_036_module_data_in[1] ;
 wire \sw_036_module_data_in[2] ;
 wire \sw_036_module_data_in[3] ;
 wire \sw_036_module_data_in[4] ;
 wire \sw_036_module_data_in[5] ;
 wire \sw_036_module_data_in[6] ;
 wire \sw_036_module_data_in[7] ;
 wire \sw_036_module_data_out[0] ;
 wire \sw_036_module_data_out[1] ;
 wire \sw_036_module_data_out[2] ;
 wire \sw_036_module_data_out[3] ;
 wire \sw_036_module_data_out[4] ;
 wire \sw_036_module_data_out[5] ;
 wire \sw_036_module_data_out[6] ;
 wire \sw_036_module_data_out[7] ;
 wire sw_036_scan_out;
 wire sw_037_clk_out;
 wire sw_037_data_out;
 wire sw_037_latch_out;
 wire \sw_037_module_data_in[0] ;
 wire \sw_037_module_data_in[1] ;
 wire \sw_037_module_data_in[2] ;
 wire \sw_037_module_data_in[3] ;
 wire \sw_037_module_data_in[4] ;
 wire \sw_037_module_data_in[5] ;
 wire \sw_037_module_data_in[6] ;
 wire \sw_037_module_data_in[7] ;
 wire \sw_037_module_data_out[0] ;
 wire \sw_037_module_data_out[1] ;
 wire \sw_037_module_data_out[2] ;
 wire \sw_037_module_data_out[3] ;
 wire \sw_037_module_data_out[4] ;
 wire \sw_037_module_data_out[5] ;
 wire \sw_037_module_data_out[6] ;
 wire \sw_037_module_data_out[7] ;
 wire sw_037_scan_out;
 wire sw_038_clk_out;
 wire sw_038_data_out;
 wire sw_038_latch_out;
 wire \sw_038_module_data_in[0] ;
 wire \sw_038_module_data_in[1] ;
 wire \sw_038_module_data_in[2] ;
 wire \sw_038_module_data_in[3] ;
 wire \sw_038_module_data_in[4] ;
 wire \sw_038_module_data_in[5] ;
 wire \sw_038_module_data_in[6] ;
 wire \sw_038_module_data_in[7] ;
 wire \sw_038_module_data_out[0] ;
 wire \sw_038_module_data_out[1] ;
 wire \sw_038_module_data_out[2] ;
 wire \sw_038_module_data_out[3] ;
 wire \sw_038_module_data_out[4] ;
 wire \sw_038_module_data_out[5] ;
 wire \sw_038_module_data_out[6] ;
 wire \sw_038_module_data_out[7] ;
 wire sw_038_scan_out;
 wire sw_039_clk_out;
 wire sw_039_data_out;
 wire sw_039_latch_out;
 wire \sw_039_module_data_in[0] ;
 wire \sw_039_module_data_in[1] ;
 wire \sw_039_module_data_in[2] ;
 wire \sw_039_module_data_in[3] ;
 wire \sw_039_module_data_in[4] ;
 wire \sw_039_module_data_in[5] ;
 wire \sw_039_module_data_in[6] ;
 wire \sw_039_module_data_in[7] ;
 wire \sw_039_module_data_out[0] ;
 wire \sw_039_module_data_out[1] ;
 wire \sw_039_module_data_out[2] ;
 wire \sw_039_module_data_out[3] ;
 wire \sw_039_module_data_out[4] ;
 wire \sw_039_module_data_out[5] ;
 wire \sw_039_module_data_out[6] ;
 wire \sw_039_module_data_out[7] ;
 wire sw_039_scan_out;
 wire sw_040_clk_out;
 wire sw_040_data_out;
 wire sw_040_latch_out;
 wire \sw_040_module_data_in[0] ;
 wire \sw_040_module_data_in[1] ;
 wire \sw_040_module_data_in[2] ;
 wire \sw_040_module_data_in[3] ;
 wire \sw_040_module_data_in[4] ;
 wire \sw_040_module_data_in[5] ;
 wire \sw_040_module_data_in[6] ;
 wire \sw_040_module_data_in[7] ;
 wire \sw_040_module_data_out[0] ;
 wire \sw_040_module_data_out[1] ;
 wire \sw_040_module_data_out[2] ;
 wire \sw_040_module_data_out[3] ;
 wire \sw_040_module_data_out[4] ;
 wire \sw_040_module_data_out[5] ;
 wire \sw_040_module_data_out[6] ;
 wire \sw_040_module_data_out[7] ;
 wire sw_040_scan_out;
 wire sw_041_clk_out;
 wire sw_041_data_out;
 wire sw_041_latch_out;
 wire \sw_041_module_data_in[0] ;
 wire \sw_041_module_data_in[1] ;
 wire \sw_041_module_data_in[2] ;
 wire \sw_041_module_data_in[3] ;
 wire \sw_041_module_data_in[4] ;
 wire \sw_041_module_data_in[5] ;
 wire \sw_041_module_data_in[6] ;
 wire \sw_041_module_data_in[7] ;
 wire \sw_041_module_data_out[0] ;
 wire \sw_041_module_data_out[1] ;
 wire \sw_041_module_data_out[2] ;
 wire \sw_041_module_data_out[3] ;
 wire \sw_041_module_data_out[4] ;
 wire \sw_041_module_data_out[5] ;
 wire \sw_041_module_data_out[6] ;
 wire \sw_041_module_data_out[7] ;
 wire sw_041_scan_out;
 wire sw_042_clk_out;
 wire sw_042_data_out;
 wire sw_042_latch_out;
 wire \sw_042_module_data_in[0] ;
 wire \sw_042_module_data_in[1] ;
 wire \sw_042_module_data_in[2] ;
 wire \sw_042_module_data_in[3] ;
 wire \sw_042_module_data_in[4] ;
 wire \sw_042_module_data_in[5] ;
 wire \sw_042_module_data_in[6] ;
 wire \sw_042_module_data_in[7] ;
 wire \sw_042_module_data_out[0] ;
 wire \sw_042_module_data_out[1] ;
 wire \sw_042_module_data_out[2] ;
 wire \sw_042_module_data_out[3] ;
 wire \sw_042_module_data_out[4] ;
 wire \sw_042_module_data_out[5] ;
 wire \sw_042_module_data_out[6] ;
 wire \sw_042_module_data_out[7] ;
 wire sw_042_scan_out;
 wire sw_043_clk_out;
 wire sw_043_data_out;
 wire sw_043_latch_out;
 wire \sw_043_module_data_in[0] ;
 wire \sw_043_module_data_in[1] ;
 wire \sw_043_module_data_in[2] ;
 wire \sw_043_module_data_in[3] ;
 wire \sw_043_module_data_in[4] ;
 wire \sw_043_module_data_in[5] ;
 wire \sw_043_module_data_in[6] ;
 wire \sw_043_module_data_in[7] ;
 wire \sw_043_module_data_out[0] ;
 wire \sw_043_module_data_out[1] ;
 wire \sw_043_module_data_out[2] ;
 wire \sw_043_module_data_out[3] ;
 wire \sw_043_module_data_out[4] ;
 wire \sw_043_module_data_out[5] ;
 wire \sw_043_module_data_out[6] ;
 wire \sw_043_module_data_out[7] ;
 wire sw_043_scan_out;
 wire sw_044_clk_out;
 wire sw_044_data_out;
 wire sw_044_latch_out;
 wire \sw_044_module_data_in[0] ;
 wire \sw_044_module_data_in[1] ;
 wire \sw_044_module_data_in[2] ;
 wire \sw_044_module_data_in[3] ;
 wire \sw_044_module_data_in[4] ;
 wire \sw_044_module_data_in[5] ;
 wire \sw_044_module_data_in[6] ;
 wire \sw_044_module_data_in[7] ;
 wire \sw_044_module_data_out[0] ;
 wire \sw_044_module_data_out[1] ;
 wire \sw_044_module_data_out[2] ;
 wire \sw_044_module_data_out[3] ;
 wire \sw_044_module_data_out[4] ;
 wire \sw_044_module_data_out[5] ;
 wire \sw_044_module_data_out[6] ;
 wire \sw_044_module_data_out[7] ;
 wire sw_044_scan_out;
 wire sw_045_clk_out;
 wire sw_045_data_out;
 wire sw_045_latch_out;
 wire \sw_045_module_data_in[0] ;
 wire \sw_045_module_data_in[1] ;
 wire \sw_045_module_data_in[2] ;
 wire \sw_045_module_data_in[3] ;
 wire \sw_045_module_data_in[4] ;
 wire \sw_045_module_data_in[5] ;
 wire \sw_045_module_data_in[6] ;
 wire \sw_045_module_data_in[7] ;
 wire \sw_045_module_data_out[0] ;
 wire \sw_045_module_data_out[1] ;
 wire \sw_045_module_data_out[2] ;
 wire \sw_045_module_data_out[3] ;
 wire \sw_045_module_data_out[4] ;
 wire \sw_045_module_data_out[5] ;
 wire \sw_045_module_data_out[6] ;
 wire \sw_045_module_data_out[7] ;
 wire sw_045_scan_out;
 wire sw_046_clk_out;
 wire sw_046_data_out;
 wire sw_046_latch_out;
 wire \sw_046_module_data_in[0] ;
 wire \sw_046_module_data_in[1] ;
 wire \sw_046_module_data_in[2] ;
 wire \sw_046_module_data_in[3] ;
 wire \sw_046_module_data_in[4] ;
 wire \sw_046_module_data_in[5] ;
 wire \sw_046_module_data_in[6] ;
 wire \sw_046_module_data_in[7] ;
 wire \sw_046_module_data_out[0] ;
 wire \sw_046_module_data_out[1] ;
 wire \sw_046_module_data_out[2] ;
 wire \sw_046_module_data_out[3] ;
 wire \sw_046_module_data_out[4] ;
 wire \sw_046_module_data_out[5] ;
 wire \sw_046_module_data_out[6] ;
 wire \sw_046_module_data_out[7] ;
 wire sw_046_scan_out;
 wire sw_047_clk_out;
 wire sw_047_data_out;
 wire sw_047_latch_out;
 wire \sw_047_module_data_in[0] ;
 wire \sw_047_module_data_in[1] ;
 wire \sw_047_module_data_in[2] ;
 wire \sw_047_module_data_in[3] ;
 wire \sw_047_module_data_in[4] ;
 wire \sw_047_module_data_in[5] ;
 wire \sw_047_module_data_in[6] ;
 wire \sw_047_module_data_in[7] ;
 wire \sw_047_module_data_out[0] ;
 wire \sw_047_module_data_out[1] ;
 wire \sw_047_module_data_out[2] ;
 wire \sw_047_module_data_out[3] ;
 wire \sw_047_module_data_out[4] ;
 wire \sw_047_module_data_out[5] ;
 wire \sw_047_module_data_out[6] ;
 wire \sw_047_module_data_out[7] ;
 wire sw_047_scan_out;
 wire sw_048_clk_out;
 wire sw_048_data_out;
 wire sw_048_latch_out;
 wire \sw_048_module_data_in[0] ;
 wire \sw_048_module_data_in[1] ;
 wire \sw_048_module_data_in[2] ;
 wire \sw_048_module_data_in[3] ;
 wire \sw_048_module_data_in[4] ;
 wire \sw_048_module_data_in[5] ;
 wire \sw_048_module_data_in[6] ;
 wire \sw_048_module_data_in[7] ;
 wire \sw_048_module_data_out[0] ;
 wire \sw_048_module_data_out[1] ;
 wire \sw_048_module_data_out[2] ;
 wire \sw_048_module_data_out[3] ;
 wire \sw_048_module_data_out[4] ;
 wire \sw_048_module_data_out[5] ;
 wire \sw_048_module_data_out[6] ;
 wire \sw_048_module_data_out[7] ;
 wire sw_048_scan_out;
 wire sw_049_clk_out;
 wire sw_049_data_out;
 wire sw_049_latch_out;
 wire \sw_049_module_data_in[0] ;
 wire \sw_049_module_data_in[1] ;
 wire \sw_049_module_data_in[2] ;
 wire \sw_049_module_data_in[3] ;
 wire \sw_049_module_data_in[4] ;
 wire \sw_049_module_data_in[5] ;
 wire \sw_049_module_data_in[6] ;
 wire \sw_049_module_data_in[7] ;
 wire \sw_049_module_data_out[0] ;
 wire \sw_049_module_data_out[1] ;
 wire \sw_049_module_data_out[2] ;
 wire \sw_049_module_data_out[3] ;
 wire \sw_049_module_data_out[4] ;
 wire \sw_049_module_data_out[5] ;
 wire \sw_049_module_data_out[6] ;
 wire \sw_049_module_data_out[7] ;
 wire sw_049_scan_out;
 wire sw_050_clk_out;
 wire sw_050_data_out;
 wire sw_050_latch_out;
 wire \sw_050_module_data_in[0] ;
 wire \sw_050_module_data_in[1] ;
 wire \sw_050_module_data_in[2] ;
 wire \sw_050_module_data_in[3] ;
 wire \sw_050_module_data_in[4] ;
 wire \sw_050_module_data_in[5] ;
 wire \sw_050_module_data_in[6] ;
 wire \sw_050_module_data_in[7] ;
 wire \sw_050_module_data_out[0] ;
 wire \sw_050_module_data_out[1] ;
 wire \sw_050_module_data_out[2] ;
 wire \sw_050_module_data_out[3] ;
 wire \sw_050_module_data_out[4] ;
 wire \sw_050_module_data_out[5] ;
 wire \sw_050_module_data_out[6] ;
 wire \sw_050_module_data_out[7] ;
 wire sw_050_scan_out;
 wire sw_051_clk_out;
 wire sw_051_data_out;
 wire sw_051_latch_out;
 wire \sw_051_module_data_in[0] ;
 wire \sw_051_module_data_in[1] ;
 wire \sw_051_module_data_in[2] ;
 wire \sw_051_module_data_in[3] ;
 wire \sw_051_module_data_in[4] ;
 wire \sw_051_module_data_in[5] ;
 wire \sw_051_module_data_in[6] ;
 wire \sw_051_module_data_in[7] ;
 wire \sw_051_module_data_out[0] ;
 wire \sw_051_module_data_out[1] ;
 wire \sw_051_module_data_out[2] ;
 wire \sw_051_module_data_out[3] ;
 wire \sw_051_module_data_out[4] ;
 wire \sw_051_module_data_out[5] ;
 wire \sw_051_module_data_out[6] ;
 wire \sw_051_module_data_out[7] ;
 wire sw_051_scan_out;
 wire sw_052_clk_out;
 wire sw_052_data_out;
 wire sw_052_latch_out;
 wire \sw_052_module_data_in[0] ;
 wire \sw_052_module_data_in[1] ;
 wire \sw_052_module_data_in[2] ;
 wire \sw_052_module_data_in[3] ;
 wire \sw_052_module_data_in[4] ;
 wire \sw_052_module_data_in[5] ;
 wire \sw_052_module_data_in[6] ;
 wire \sw_052_module_data_in[7] ;
 wire \sw_052_module_data_out[0] ;
 wire \sw_052_module_data_out[1] ;
 wire \sw_052_module_data_out[2] ;
 wire \sw_052_module_data_out[3] ;
 wire \sw_052_module_data_out[4] ;
 wire \sw_052_module_data_out[5] ;
 wire \sw_052_module_data_out[6] ;
 wire \sw_052_module_data_out[7] ;
 wire sw_052_scan_out;
 wire sw_053_clk_out;
 wire sw_053_data_out;
 wire sw_053_latch_out;
 wire \sw_053_module_data_in[0] ;
 wire \sw_053_module_data_in[1] ;
 wire \sw_053_module_data_in[2] ;
 wire \sw_053_module_data_in[3] ;
 wire \sw_053_module_data_in[4] ;
 wire \sw_053_module_data_in[5] ;
 wire \sw_053_module_data_in[6] ;
 wire \sw_053_module_data_in[7] ;
 wire \sw_053_module_data_out[0] ;
 wire \sw_053_module_data_out[1] ;
 wire \sw_053_module_data_out[2] ;
 wire \sw_053_module_data_out[3] ;
 wire \sw_053_module_data_out[4] ;
 wire \sw_053_module_data_out[5] ;
 wire \sw_053_module_data_out[6] ;
 wire \sw_053_module_data_out[7] ;
 wire sw_053_scan_out;
 wire sw_054_clk_out;
 wire sw_054_data_out;
 wire sw_054_latch_out;
 wire \sw_054_module_data_in[0] ;
 wire \sw_054_module_data_in[1] ;
 wire \sw_054_module_data_in[2] ;
 wire \sw_054_module_data_in[3] ;
 wire \sw_054_module_data_in[4] ;
 wire \sw_054_module_data_in[5] ;
 wire \sw_054_module_data_in[6] ;
 wire \sw_054_module_data_in[7] ;
 wire \sw_054_module_data_out[0] ;
 wire \sw_054_module_data_out[1] ;
 wire \sw_054_module_data_out[2] ;
 wire \sw_054_module_data_out[3] ;
 wire \sw_054_module_data_out[4] ;
 wire \sw_054_module_data_out[5] ;
 wire \sw_054_module_data_out[6] ;
 wire \sw_054_module_data_out[7] ;
 wire sw_054_scan_out;
 wire sw_055_clk_out;
 wire sw_055_data_out;
 wire sw_055_latch_out;
 wire \sw_055_module_data_in[0] ;
 wire \sw_055_module_data_in[1] ;
 wire \sw_055_module_data_in[2] ;
 wire \sw_055_module_data_in[3] ;
 wire \sw_055_module_data_in[4] ;
 wire \sw_055_module_data_in[5] ;
 wire \sw_055_module_data_in[6] ;
 wire \sw_055_module_data_in[7] ;
 wire \sw_055_module_data_out[0] ;
 wire \sw_055_module_data_out[1] ;
 wire \sw_055_module_data_out[2] ;
 wire \sw_055_module_data_out[3] ;
 wire \sw_055_module_data_out[4] ;
 wire \sw_055_module_data_out[5] ;
 wire \sw_055_module_data_out[6] ;
 wire \sw_055_module_data_out[7] ;
 wire sw_055_scan_out;
 wire sw_056_clk_out;
 wire sw_056_data_out;
 wire sw_056_latch_out;
 wire \sw_056_module_data_in[0] ;
 wire \sw_056_module_data_in[1] ;
 wire \sw_056_module_data_in[2] ;
 wire \sw_056_module_data_in[3] ;
 wire \sw_056_module_data_in[4] ;
 wire \sw_056_module_data_in[5] ;
 wire \sw_056_module_data_in[6] ;
 wire \sw_056_module_data_in[7] ;
 wire \sw_056_module_data_out[0] ;
 wire \sw_056_module_data_out[1] ;
 wire \sw_056_module_data_out[2] ;
 wire \sw_056_module_data_out[3] ;
 wire \sw_056_module_data_out[4] ;
 wire \sw_056_module_data_out[5] ;
 wire \sw_056_module_data_out[6] ;
 wire \sw_056_module_data_out[7] ;
 wire sw_056_scan_out;
 wire sw_057_clk_out;
 wire sw_057_data_out;
 wire sw_057_latch_out;
 wire \sw_057_module_data_in[0] ;
 wire \sw_057_module_data_in[1] ;
 wire \sw_057_module_data_in[2] ;
 wire \sw_057_module_data_in[3] ;
 wire \sw_057_module_data_in[4] ;
 wire \sw_057_module_data_in[5] ;
 wire \sw_057_module_data_in[6] ;
 wire \sw_057_module_data_in[7] ;
 wire \sw_057_module_data_out[0] ;
 wire \sw_057_module_data_out[1] ;
 wire \sw_057_module_data_out[2] ;
 wire \sw_057_module_data_out[3] ;
 wire \sw_057_module_data_out[4] ;
 wire \sw_057_module_data_out[5] ;
 wire \sw_057_module_data_out[6] ;
 wire \sw_057_module_data_out[7] ;
 wire sw_057_scan_out;
 wire sw_058_clk_out;
 wire sw_058_data_out;
 wire sw_058_latch_out;
 wire \sw_058_module_data_in[0] ;
 wire \sw_058_module_data_in[1] ;
 wire \sw_058_module_data_in[2] ;
 wire \sw_058_module_data_in[3] ;
 wire \sw_058_module_data_in[4] ;
 wire \sw_058_module_data_in[5] ;
 wire \sw_058_module_data_in[6] ;
 wire \sw_058_module_data_in[7] ;
 wire \sw_058_module_data_out[0] ;
 wire \sw_058_module_data_out[1] ;
 wire \sw_058_module_data_out[2] ;
 wire \sw_058_module_data_out[3] ;
 wire \sw_058_module_data_out[4] ;
 wire \sw_058_module_data_out[5] ;
 wire \sw_058_module_data_out[6] ;
 wire \sw_058_module_data_out[7] ;
 wire sw_058_scan_out;
 wire sw_059_clk_out;
 wire sw_059_data_out;
 wire sw_059_latch_out;
 wire \sw_059_module_data_in[0] ;
 wire \sw_059_module_data_in[1] ;
 wire \sw_059_module_data_in[2] ;
 wire \sw_059_module_data_in[3] ;
 wire \sw_059_module_data_in[4] ;
 wire \sw_059_module_data_in[5] ;
 wire \sw_059_module_data_in[6] ;
 wire \sw_059_module_data_in[7] ;
 wire \sw_059_module_data_out[0] ;
 wire \sw_059_module_data_out[1] ;
 wire \sw_059_module_data_out[2] ;
 wire \sw_059_module_data_out[3] ;
 wire \sw_059_module_data_out[4] ;
 wire \sw_059_module_data_out[5] ;
 wire \sw_059_module_data_out[6] ;
 wire \sw_059_module_data_out[7] ;
 wire sw_059_scan_out;
 wire sw_060_clk_out;
 wire sw_060_data_out;
 wire sw_060_latch_out;
 wire \sw_060_module_data_in[0] ;
 wire \sw_060_module_data_in[1] ;
 wire \sw_060_module_data_in[2] ;
 wire \sw_060_module_data_in[3] ;
 wire \sw_060_module_data_in[4] ;
 wire \sw_060_module_data_in[5] ;
 wire \sw_060_module_data_in[6] ;
 wire \sw_060_module_data_in[7] ;
 wire \sw_060_module_data_out[0] ;
 wire \sw_060_module_data_out[1] ;
 wire \sw_060_module_data_out[2] ;
 wire \sw_060_module_data_out[3] ;
 wire \sw_060_module_data_out[4] ;
 wire \sw_060_module_data_out[5] ;
 wire \sw_060_module_data_out[6] ;
 wire \sw_060_module_data_out[7] ;
 wire sw_060_scan_out;
 wire sw_061_clk_out;
 wire sw_061_data_out;
 wire sw_061_latch_out;
 wire \sw_061_module_data_in[0] ;
 wire \sw_061_module_data_in[1] ;
 wire \sw_061_module_data_in[2] ;
 wire \sw_061_module_data_in[3] ;
 wire \sw_061_module_data_in[4] ;
 wire \sw_061_module_data_in[5] ;
 wire \sw_061_module_data_in[6] ;
 wire \sw_061_module_data_in[7] ;
 wire \sw_061_module_data_out[0] ;
 wire \sw_061_module_data_out[1] ;
 wire \sw_061_module_data_out[2] ;
 wire \sw_061_module_data_out[3] ;
 wire \sw_061_module_data_out[4] ;
 wire \sw_061_module_data_out[5] ;
 wire \sw_061_module_data_out[6] ;
 wire \sw_061_module_data_out[7] ;
 wire sw_061_scan_out;
 wire sw_062_clk_out;
 wire sw_062_data_out;
 wire sw_062_latch_out;
 wire \sw_062_module_data_in[0] ;
 wire \sw_062_module_data_in[1] ;
 wire \sw_062_module_data_in[2] ;
 wire \sw_062_module_data_in[3] ;
 wire \sw_062_module_data_in[4] ;
 wire \sw_062_module_data_in[5] ;
 wire \sw_062_module_data_in[6] ;
 wire \sw_062_module_data_in[7] ;
 wire \sw_062_module_data_out[0] ;
 wire \sw_062_module_data_out[1] ;
 wire \sw_062_module_data_out[2] ;
 wire \sw_062_module_data_out[3] ;
 wire \sw_062_module_data_out[4] ;
 wire \sw_062_module_data_out[5] ;
 wire \sw_062_module_data_out[6] ;
 wire \sw_062_module_data_out[7] ;
 wire sw_062_scan_out;
 wire sw_063_clk_out;
 wire sw_063_data_out;
 wire sw_063_latch_out;
 wire \sw_063_module_data_in[0] ;
 wire \sw_063_module_data_in[1] ;
 wire \sw_063_module_data_in[2] ;
 wire \sw_063_module_data_in[3] ;
 wire \sw_063_module_data_in[4] ;
 wire \sw_063_module_data_in[5] ;
 wire \sw_063_module_data_in[6] ;
 wire \sw_063_module_data_in[7] ;
 wire \sw_063_module_data_out[0] ;
 wire \sw_063_module_data_out[1] ;
 wire \sw_063_module_data_out[2] ;
 wire \sw_063_module_data_out[3] ;
 wire \sw_063_module_data_out[4] ;
 wire \sw_063_module_data_out[5] ;
 wire \sw_063_module_data_out[6] ;
 wire \sw_063_module_data_out[7] ;
 wire sw_063_scan_out;
 wire sw_064_clk_out;
 wire sw_064_data_out;
 wire sw_064_latch_out;
 wire \sw_064_module_data_in[0] ;
 wire \sw_064_module_data_in[1] ;
 wire \sw_064_module_data_in[2] ;
 wire \sw_064_module_data_in[3] ;
 wire \sw_064_module_data_in[4] ;
 wire \sw_064_module_data_in[5] ;
 wire \sw_064_module_data_in[6] ;
 wire \sw_064_module_data_in[7] ;
 wire \sw_064_module_data_out[0] ;
 wire \sw_064_module_data_out[1] ;
 wire \sw_064_module_data_out[2] ;
 wire \sw_064_module_data_out[3] ;
 wire \sw_064_module_data_out[4] ;
 wire \sw_064_module_data_out[5] ;
 wire \sw_064_module_data_out[6] ;
 wire \sw_064_module_data_out[7] ;
 wire sw_064_scan_out;
 wire sw_065_clk_out;
 wire sw_065_data_out;
 wire sw_065_latch_out;
 wire \sw_065_module_data_in[0] ;
 wire \sw_065_module_data_in[1] ;
 wire \sw_065_module_data_in[2] ;
 wire \sw_065_module_data_in[3] ;
 wire \sw_065_module_data_in[4] ;
 wire \sw_065_module_data_in[5] ;
 wire \sw_065_module_data_in[6] ;
 wire \sw_065_module_data_in[7] ;
 wire \sw_065_module_data_out[0] ;
 wire \sw_065_module_data_out[1] ;
 wire \sw_065_module_data_out[2] ;
 wire \sw_065_module_data_out[3] ;
 wire \sw_065_module_data_out[4] ;
 wire \sw_065_module_data_out[5] ;
 wire \sw_065_module_data_out[6] ;
 wire \sw_065_module_data_out[7] ;
 wire sw_065_scan_out;
 wire sw_066_clk_out;
 wire sw_066_data_out;
 wire sw_066_latch_out;
 wire \sw_066_module_data_in[0] ;
 wire \sw_066_module_data_in[1] ;
 wire \sw_066_module_data_in[2] ;
 wire \sw_066_module_data_in[3] ;
 wire \sw_066_module_data_in[4] ;
 wire \sw_066_module_data_in[5] ;
 wire \sw_066_module_data_in[6] ;
 wire \sw_066_module_data_in[7] ;
 wire \sw_066_module_data_out[0] ;
 wire \sw_066_module_data_out[1] ;
 wire \sw_066_module_data_out[2] ;
 wire \sw_066_module_data_out[3] ;
 wire \sw_066_module_data_out[4] ;
 wire \sw_066_module_data_out[5] ;
 wire \sw_066_module_data_out[6] ;
 wire \sw_066_module_data_out[7] ;
 wire sw_066_scan_out;
 wire sw_067_clk_out;
 wire sw_067_data_out;
 wire sw_067_latch_out;
 wire \sw_067_module_data_in[0] ;
 wire \sw_067_module_data_in[1] ;
 wire \sw_067_module_data_in[2] ;
 wire \sw_067_module_data_in[3] ;
 wire \sw_067_module_data_in[4] ;
 wire \sw_067_module_data_in[5] ;
 wire \sw_067_module_data_in[6] ;
 wire \sw_067_module_data_in[7] ;
 wire \sw_067_module_data_out[0] ;
 wire \sw_067_module_data_out[1] ;
 wire \sw_067_module_data_out[2] ;
 wire \sw_067_module_data_out[3] ;
 wire \sw_067_module_data_out[4] ;
 wire \sw_067_module_data_out[5] ;
 wire \sw_067_module_data_out[6] ;
 wire \sw_067_module_data_out[7] ;
 wire sw_067_scan_out;
 wire sw_068_clk_out;
 wire sw_068_data_out;
 wire sw_068_latch_out;
 wire \sw_068_module_data_in[0] ;
 wire \sw_068_module_data_in[1] ;
 wire \sw_068_module_data_in[2] ;
 wire \sw_068_module_data_in[3] ;
 wire \sw_068_module_data_in[4] ;
 wire \sw_068_module_data_in[5] ;
 wire \sw_068_module_data_in[6] ;
 wire \sw_068_module_data_in[7] ;
 wire \sw_068_module_data_out[0] ;
 wire \sw_068_module_data_out[1] ;
 wire \sw_068_module_data_out[2] ;
 wire \sw_068_module_data_out[3] ;
 wire \sw_068_module_data_out[4] ;
 wire \sw_068_module_data_out[5] ;
 wire \sw_068_module_data_out[6] ;
 wire \sw_068_module_data_out[7] ;
 wire sw_068_scan_out;
 wire sw_069_clk_out;
 wire sw_069_data_out;
 wire sw_069_latch_out;
 wire \sw_069_module_data_in[0] ;
 wire \sw_069_module_data_in[1] ;
 wire \sw_069_module_data_in[2] ;
 wire \sw_069_module_data_in[3] ;
 wire \sw_069_module_data_in[4] ;
 wire \sw_069_module_data_in[5] ;
 wire \sw_069_module_data_in[6] ;
 wire \sw_069_module_data_in[7] ;
 wire \sw_069_module_data_out[0] ;
 wire \sw_069_module_data_out[1] ;
 wire \sw_069_module_data_out[2] ;
 wire \sw_069_module_data_out[3] ;
 wire \sw_069_module_data_out[4] ;
 wire \sw_069_module_data_out[5] ;
 wire \sw_069_module_data_out[6] ;
 wire \sw_069_module_data_out[7] ;
 wire sw_069_scan_out;
 wire sw_070_clk_out;
 wire sw_070_data_out;
 wire sw_070_latch_out;
 wire \sw_070_module_data_in[0] ;
 wire \sw_070_module_data_in[1] ;
 wire \sw_070_module_data_in[2] ;
 wire \sw_070_module_data_in[3] ;
 wire \sw_070_module_data_in[4] ;
 wire \sw_070_module_data_in[5] ;
 wire \sw_070_module_data_in[6] ;
 wire \sw_070_module_data_in[7] ;
 wire \sw_070_module_data_out[0] ;
 wire \sw_070_module_data_out[1] ;
 wire \sw_070_module_data_out[2] ;
 wire \sw_070_module_data_out[3] ;
 wire \sw_070_module_data_out[4] ;
 wire \sw_070_module_data_out[5] ;
 wire \sw_070_module_data_out[6] ;
 wire \sw_070_module_data_out[7] ;
 wire sw_070_scan_out;
 wire sw_071_clk_out;
 wire sw_071_data_out;
 wire sw_071_latch_out;
 wire \sw_071_module_data_in[0] ;
 wire \sw_071_module_data_in[1] ;
 wire \sw_071_module_data_in[2] ;
 wire \sw_071_module_data_in[3] ;
 wire \sw_071_module_data_in[4] ;
 wire \sw_071_module_data_in[5] ;
 wire \sw_071_module_data_in[6] ;
 wire \sw_071_module_data_in[7] ;
 wire \sw_071_module_data_out[0] ;
 wire \sw_071_module_data_out[1] ;
 wire \sw_071_module_data_out[2] ;
 wire \sw_071_module_data_out[3] ;
 wire \sw_071_module_data_out[4] ;
 wire \sw_071_module_data_out[5] ;
 wire \sw_071_module_data_out[6] ;
 wire \sw_071_module_data_out[7] ;
 wire sw_071_scan_out;
 wire sw_072_clk_out;
 wire sw_072_data_out;
 wire sw_072_latch_out;
 wire \sw_072_module_data_in[0] ;
 wire \sw_072_module_data_in[1] ;
 wire \sw_072_module_data_in[2] ;
 wire \sw_072_module_data_in[3] ;
 wire \sw_072_module_data_in[4] ;
 wire \sw_072_module_data_in[5] ;
 wire \sw_072_module_data_in[6] ;
 wire \sw_072_module_data_in[7] ;
 wire \sw_072_module_data_out[0] ;
 wire \sw_072_module_data_out[1] ;
 wire \sw_072_module_data_out[2] ;
 wire \sw_072_module_data_out[3] ;
 wire \sw_072_module_data_out[4] ;
 wire \sw_072_module_data_out[5] ;
 wire \sw_072_module_data_out[6] ;
 wire \sw_072_module_data_out[7] ;
 wire sw_072_scan_out;
 wire sw_073_clk_out;
 wire sw_073_data_out;
 wire sw_073_latch_out;
 wire \sw_073_module_data_in[0] ;
 wire \sw_073_module_data_in[1] ;
 wire \sw_073_module_data_in[2] ;
 wire \sw_073_module_data_in[3] ;
 wire \sw_073_module_data_in[4] ;
 wire \sw_073_module_data_in[5] ;
 wire \sw_073_module_data_in[6] ;
 wire \sw_073_module_data_in[7] ;
 wire \sw_073_module_data_out[0] ;
 wire \sw_073_module_data_out[1] ;
 wire \sw_073_module_data_out[2] ;
 wire \sw_073_module_data_out[3] ;
 wire \sw_073_module_data_out[4] ;
 wire \sw_073_module_data_out[5] ;
 wire \sw_073_module_data_out[6] ;
 wire \sw_073_module_data_out[7] ;
 wire sw_073_scan_out;
 wire sw_074_clk_out;
 wire sw_074_data_out;
 wire sw_074_latch_out;
 wire \sw_074_module_data_in[0] ;
 wire \sw_074_module_data_in[1] ;
 wire \sw_074_module_data_in[2] ;
 wire \sw_074_module_data_in[3] ;
 wire \sw_074_module_data_in[4] ;
 wire \sw_074_module_data_in[5] ;
 wire \sw_074_module_data_in[6] ;
 wire \sw_074_module_data_in[7] ;
 wire \sw_074_module_data_out[0] ;
 wire \sw_074_module_data_out[1] ;
 wire \sw_074_module_data_out[2] ;
 wire \sw_074_module_data_out[3] ;
 wire \sw_074_module_data_out[4] ;
 wire \sw_074_module_data_out[5] ;
 wire \sw_074_module_data_out[6] ;
 wire \sw_074_module_data_out[7] ;
 wire sw_074_scan_out;
 wire sw_075_clk_out;
 wire sw_075_data_out;
 wire sw_075_latch_out;
 wire \sw_075_module_data_in[0] ;
 wire \sw_075_module_data_in[1] ;
 wire \sw_075_module_data_in[2] ;
 wire \sw_075_module_data_in[3] ;
 wire \sw_075_module_data_in[4] ;
 wire \sw_075_module_data_in[5] ;
 wire \sw_075_module_data_in[6] ;
 wire \sw_075_module_data_in[7] ;
 wire \sw_075_module_data_out[0] ;
 wire \sw_075_module_data_out[1] ;
 wire \sw_075_module_data_out[2] ;
 wire \sw_075_module_data_out[3] ;
 wire \sw_075_module_data_out[4] ;
 wire \sw_075_module_data_out[5] ;
 wire \sw_075_module_data_out[6] ;
 wire \sw_075_module_data_out[7] ;
 wire sw_075_scan_out;
 wire sw_076_clk_out;
 wire sw_076_data_out;
 wire sw_076_latch_out;
 wire \sw_076_module_data_in[0] ;
 wire \sw_076_module_data_in[1] ;
 wire \sw_076_module_data_in[2] ;
 wire \sw_076_module_data_in[3] ;
 wire \sw_076_module_data_in[4] ;
 wire \sw_076_module_data_in[5] ;
 wire \sw_076_module_data_in[6] ;
 wire \sw_076_module_data_in[7] ;
 wire \sw_076_module_data_out[0] ;
 wire \sw_076_module_data_out[1] ;
 wire \sw_076_module_data_out[2] ;
 wire \sw_076_module_data_out[3] ;
 wire \sw_076_module_data_out[4] ;
 wire \sw_076_module_data_out[5] ;
 wire \sw_076_module_data_out[6] ;
 wire \sw_076_module_data_out[7] ;
 wire sw_076_scan_out;
 wire sw_077_clk_out;
 wire sw_077_data_out;
 wire sw_077_latch_out;
 wire \sw_077_module_data_in[0] ;
 wire \sw_077_module_data_in[1] ;
 wire \sw_077_module_data_in[2] ;
 wire \sw_077_module_data_in[3] ;
 wire \sw_077_module_data_in[4] ;
 wire \sw_077_module_data_in[5] ;
 wire \sw_077_module_data_in[6] ;
 wire \sw_077_module_data_in[7] ;
 wire \sw_077_module_data_out[0] ;
 wire \sw_077_module_data_out[1] ;
 wire \sw_077_module_data_out[2] ;
 wire \sw_077_module_data_out[3] ;
 wire \sw_077_module_data_out[4] ;
 wire \sw_077_module_data_out[5] ;
 wire \sw_077_module_data_out[6] ;
 wire \sw_077_module_data_out[7] ;
 wire sw_077_scan_out;
 wire sw_078_clk_out;
 wire sw_078_data_out;
 wire sw_078_latch_out;
 wire \sw_078_module_data_in[0] ;
 wire \sw_078_module_data_in[1] ;
 wire \sw_078_module_data_in[2] ;
 wire \sw_078_module_data_in[3] ;
 wire \sw_078_module_data_in[4] ;
 wire \sw_078_module_data_in[5] ;
 wire \sw_078_module_data_in[6] ;
 wire \sw_078_module_data_in[7] ;
 wire \sw_078_module_data_out[0] ;
 wire \sw_078_module_data_out[1] ;
 wire \sw_078_module_data_out[2] ;
 wire \sw_078_module_data_out[3] ;
 wire \sw_078_module_data_out[4] ;
 wire \sw_078_module_data_out[5] ;
 wire \sw_078_module_data_out[6] ;
 wire \sw_078_module_data_out[7] ;
 wire sw_078_scan_out;
 wire sw_079_clk_out;
 wire sw_079_data_out;
 wire sw_079_latch_out;
 wire \sw_079_module_data_in[0] ;
 wire \sw_079_module_data_in[1] ;
 wire \sw_079_module_data_in[2] ;
 wire \sw_079_module_data_in[3] ;
 wire \sw_079_module_data_in[4] ;
 wire \sw_079_module_data_in[5] ;
 wire \sw_079_module_data_in[6] ;
 wire \sw_079_module_data_in[7] ;
 wire \sw_079_module_data_out[0] ;
 wire \sw_079_module_data_out[1] ;
 wire \sw_079_module_data_out[2] ;
 wire \sw_079_module_data_out[3] ;
 wire \sw_079_module_data_out[4] ;
 wire \sw_079_module_data_out[5] ;
 wire \sw_079_module_data_out[6] ;
 wire \sw_079_module_data_out[7] ;
 wire sw_079_scan_out;
 wire sw_080_clk_out;
 wire sw_080_data_out;
 wire sw_080_latch_out;
 wire \sw_080_module_data_in[0] ;
 wire \sw_080_module_data_in[1] ;
 wire \sw_080_module_data_in[2] ;
 wire \sw_080_module_data_in[3] ;
 wire \sw_080_module_data_in[4] ;
 wire \sw_080_module_data_in[5] ;
 wire \sw_080_module_data_in[6] ;
 wire \sw_080_module_data_in[7] ;
 wire \sw_080_module_data_out[0] ;
 wire \sw_080_module_data_out[1] ;
 wire \sw_080_module_data_out[2] ;
 wire \sw_080_module_data_out[3] ;
 wire \sw_080_module_data_out[4] ;
 wire \sw_080_module_data_out[5] ;
 wire \sw_080_module_data_out[6] ;
 wire \sw_080_module_data_out[7] ;
 wire sw_080_scan_out;
 wire sw_081_clk_out;
 wire sw_081_data_out;
 wire sw_081_latch_out;
 wire \sw_081_module_data_in[0] ;
 wire \sw_081_module_data_in[1] ;
 wire \sw_081_module_data_in[2] ;
 wire \sw_081_module_data_in[3] ;
 wire \sw_081_module_data_in[4] ;
 wire \sw_081_module_data_in[5] ;
 wire \sw_081_module_data_in[6] ;
 wire \sw_081_module_data_in[7] ;
 wire \sw_081_module_data_out[0] ;
 wire \sw_081_module_data_out[1] ;
 wire \sw_081_module_data_out[2] ;
 wire \sw_081_module_data_out[3] ;
 wire \sw_081_module_data_out[4] ;
 wire \sw_081_module_data_out[5] ;
 wire \sw_081_module_data_out[6] ;
 wire \sw_081_module_data_out[7] ;
 wire sw_081_scan_out;
 wire sw_082_clk_out;
 wire sw_082_data_out;
 wire sw_082_latch_out;
 wire \sw_082_module_data_in[0] ;
 wire \sw_082_module_data_in[1] ;
 wire \sw_082_module_data_in[2] ;
 wire \sw_082_module_data_in[3] ;
 wire \sw_082_module_data_in[4] ;
 wire \sw_082_module_data_in[5] ;
 wire \sw_082_module_data_in[6] ;
 wire \sw_082_module_data_in[7] ;
 wire \sw_082_module_data_out[0] ;
 wire \sw_082_module_data_out[1] ;
 wire \sw_082_module_data_out[2] ;
 wire \sw_082_module_data_out[3] ;
 wire \sw_082_module_data_out[4] ;
 wire \sw_082_module_data_out[5] ;
 wire \sw_082_module_data_out[6] ;
 wire \sw_082_module_data_out[7] ;
 wire sw_082_scan_out;
 wire sw_083_clk_out;
 wire sw_083_data_out;
 wire sw_083_latch_out;
 wire \sw_083_module_data_in[0] ;
 wire \sw_083_module_data_in[1] ;
 wire \sw_083_module_data_in[2] ;
 wire \sw_083_module_data_in[3] ;
 wire \sw_083_module_data_in[4] ;
 wire \sw_083_module_data_in[5] ;
 wire \sw_083_module_data_in[6] ;
 wire \sw_083_module_data_in[7] ;
 wire \sw_083_module_data_out[0] ;
 wire \sw_083_module_data_out[1] ;
 wire \sw_083_module_data_out[2] ;
 wire \sw_083_module_data_out[3] ;
 wire \sw_083_module_data_out[4] ;
 wire \sw_083_module_data_out[5] ;
 wire \sw_083_module_data_out[6] ;
 wire \sw_083_module_data_out[7] ;
 wire sw_083_scan_out;
 wire sw_084_clk_out;
 wire sw_084_data_out;
 wire sw_084_latch_out;
 wire \sw_084_module_data_in[0] ;
 wire \sw_084_module_data_in[1] ;
 wire \sw_084_module_data_in[2] ;
 wire \sw_084_module_data_in[3] ;
 wire \sw_084_module_data_in[4] ;
 wire \sw_084_module_data_in[5] ;
 wire \sw_084_module_data_in[6] ;
 wire \sw_084_module_data_in[7] ;
 wire \sw_084_module_data_out[0] ;
 wire \sw_084_module_data_out[1] ;
 wire \sw_084_module_data_out[2] ;
 wire \sw_084_module_data_out[3] ;
 wire \sw_084_module_data_out[4] ;
 wire \sw_084_module_data_out[5] ;
 wire \sw_084_module_data_out[6] ;
 wire \sw_084_module_data_out[7] ;
 wire sw_084_scan_out;
 wire sw_085_clk_out;
 wire sw_085_data_out;
 wire sw_085_latch_out;
 wire \sw_085_module_data_in[0] ;
 wire \sw_085_module_data_in[1] ;
 wire \sw_085_module_data_in[2] ;
 wire \sw_085_module_data_in[3] ;
 wire \sw_085_module_data_in[4] ;
 wire \sw_085_module_data_in[5] ;
 wire \sw_085_module_data_in[6] ;
 wire \sw_085_module_data_in[7] ;
 wire \sw_085_module_data_out[0] ;
 wire \sw_085_module_data_out[1] ;
 wire \sw_085_module_data_out[2] ;
 wire \sw_085_module_data_out[3] ;
 wire \sw_085_module_data_out[4] ;
 wire \sw_085_module_data_out[5] ;
 wire \sw_085_module_data_out[6] ;
 wire \sw_085_module_data_out[7] ;
 wire sw_085_scan_out;
 wire sw_086_clk_out;
 wire sw_086_data_out;
 wire sw_086_latch_out;
 wire \sw_086_module_data_in[0] ;
 wire \sw_086_module_data_in[1] ;
 wire \sw_086_module_data_in[2] ;
 wire \sw_086_module_data_in[3] ;
 wire \sw_086_module_data_in[4] ;
 wire \sw_086_module_data_in[5] ;
 wire \sw_086_module_data_in[6] ;
 wire \sw_086_module_data_in[7] ;
 wire \sw_086_module_data_out[0] ;
 wire \sw_086_module_data_out[1] ;
 wire \sw_086_module_data_out[2] ;
 wire \sw_086_module_data_out[3] ;
 wire \sw_086_module_data_out[4] ;
 wire \sw_086_module_data_out[5] ;
 wire \sw_086_module_data_out[6] ;
 wire \sw_086_module_data_out[7] ;
 wire sw_086_scan_out;
 wire sw_087_clk_out;
 wire sw_087_data_out;
 wire sw_087_latch_out;
 wire \sw_087_module_data_in[0] ;
 wire \sw_087_module_data_in[1] ;
 wire \sw_087_module_data_in[2] ;
 wire \sw_087_module_data_in[3] ;
 wire \sw_087_module_data_in[4] ;
 wire \sw_087_module_data_in[5] ;
 wire \sw_087_module_data_in[6] ;
 wire \sw_087_module_data_in[7] ;
 wire \sw_087_module_data_out[0] ;
 wire \sw_087_module_data_out[1] ;
 wire \sw_087_module_data_out[2] ;
 wire \sw_087_module_data_out[3] ;
 wire \sw_087_module_data_out[4] ;
 wire \sw_087_module_data_out[5] ;
 wire \sw_087_module_data_out[6] ;
 wire \sw_087_module_data_out[7] ;
 wire sw_087_scan_out;
 wire sw_088_clk_out;
 wire sw_088_data_out;
 wire sw_088_latch_out;
 wire \sw_088_module_data_in[0] ;
 wire \sw_088_module_data_in[1] ;
 wire \sw_088_module_data_in[2] ;
 wire \sw_088_module_data_in[3] ;
 wire \sw_088_module_data_in[4] ;
 wire \sw_088_module_data_in[5] ;
 wire \sw_088_module_data_in[6] ;
 wire \sw_088_module_data_in[7] ;
 wire \sw_088_module_data_out[0] ;
 wire \sw_088_module_data_out[1] ;
 wire \sw_088_module_data_out[2] ;
 wire \sw_088_module_data_out[3] ;
 wire \sw_088_module_data_out[4] ;
 wire \sw_088_module_data_out[5] ;
 wire \sw_088_module_data_out[6] ;
 wire \sw_088_module_data_out[7] ;
 wire sw_088_scan_out;
 wire sw_089_clk_out;
 wire sw_089_data_out;
 wire sw_089_latch_out;
 wire \sw_089_module_data_in[0] ;
 wire \sw_089_module_data_in[1] ;
 wire \sw_089_module_data_in[2] ;
 wire \sw_089_module_data_in[3] ;
 wire \sw_089_module_data_in[4] ;
 wire \sw_089_module_data_in[5] ;
 wire \sw_089_module_data_in[6] ;
 wire \sw_089_module_data_in[7] ;
 wire \sw_089_module_data_out[0] ;
 wire \sw_089_module_data_out[1] ;
 wire \sw_089_module_data_out[2] ;
 wire \sw_089_module_data_out[3] ;
 wire \sw_089_module_data_out[4] ;
 wire \sw_089_module_data_out[5] ;
 wire \sw_089_module_data_out[6] ;
 wire \sw_089_module_data_out[7] ;
 wire sw_089_scan_out;
 wire sw_090_clk_out;
 wire sw_090_data_out;
 wire sw_090_latch_out;
 wire \sw_090_module_data_in[0] ;
 wire \sw_090_module_data_in[1] ;
 wire \sw_090_module_data_in[2] ;
 wire \sw_090_module_data_in[3] ;
 wire \sw_090_module_data_in[4] ;
 wire \sw_090_module_data_in[5] ;
 wire \sw_090_module_data_in[6] ;
 wire \sw_090_module_data_in[7] ;
 wire \sw_090_module_data_out[0] ;
 wire \sw_090_module_data_out[1] ;
 wire \sw_090_module_data_out[2] ;
 wire \sw_090_module_data_out[3] ;
 wire \sw_090_module_data_out[4] ;
 wire \sw_090_module_data_out[5] ;
 wire \sw_090_module_data_out[6] ;
 wire \sw_090_module_data_out[7] ;
 wire sw_090_scan_out;
 wire sw_091_clk_out;
 wire sw_091_data_out;
 wire sw_091_latch_out;
 wire \sw_091_module_data_in[0] ;
 wire \sw_091_module_data_in[1] ;
 wire \sw_091_module_data_in[2] ;
 wire \sw_091_module_data_in[3] ;
 wire \sw_091_module_data_in[4] ;
 wire \sw_091_module_data_in[5] ;
 wire \sw_091_module_data_in[6] ;
 wire \sw_091_module_data_in[7] ;
 wire \sw_091_module_data_out[0] ;
 wire \sw_091_module_data_out[1] ;
 wire \sw_091_module_data_out[2] ;
 wire \sw_091_module_data_out[3] ;
 wire \sw_091_module_data_out[4] ;
 wire \sw_091_module_data_out[5] ;
 wire \sw_091_module_data_out[6] ;
 wire \sw_091_module_data_out[7] ;
 wire sw_091_scan_out;
 wire sw_092_clk_out;
 wire sw_092_data_out;
 wire sw_092_latch_out;
 wire \sw_092_module_data_in[0] ;
 wire \sw_092_module_data_in[1] ;
 wire \sw_092_module_data_in[2] ;
 wire \sw_092_module_data_in[3] ;
 wire \sw_092_module_data_in[4] ;
 wire \sw_092_module_data_in[5] ;
 wire \sw_092_module_data_in[6] ;
 wire \sw_092_module_data_in[7] ;
 wire \sw_092_module_data_out[0] ;
 wire \sw_092_module_data_out[1] ;
 wire \sw_092_module_data_out[2] ;
 wire \sw_092_module_data_out[3] ;
 wire \sw_092_module_data_out[4] ;
 wire \sw_092_module_data_out[5] ;
 wire \sw_092_module_data_out[6] ;
 wire \sw_092_module_data_out[7] ;
 wire sw_092_scan_out;
 wire sw_093_clk_out;
 wire sw_093_data_out;
 wire sw_093_latch_out;
 wire \sw_093_module_data_in[0] ;
 wire \sw_093_module_data_in[1] ;
 wire \sw_093_module_data_in[2] ;
 wire \sw_093_module_data_in[3] ;
 wire \sw_093_module_data_in[4] ;
 wire \sw_093_module_data_in[5] ;
 wire \sw_093_module_data_in[6] ;
 wire \sw_093_module_data_in[7] ;
 wire \sw_093_module_data_out[0] ;
 wire \sw_093_module_data_out[1] ;
 wire \sw_093_module_data_out[2] ;
 wire \sw_093_module_data_out[3] ;
 wire \sw_093_module_data_out[4] ;
 wire \sw_093_module_data_out[5] ;
 wire \sw_093_module_data_out[6] ;
 wire \sw_093_module_data_out[7] ;
 wire sw_093_scan_out;
 wire sw_094_clk_out;
 wire sw_094_data_out;
 wire sw_094_latch_out;
 wire \sw_094_module_data_in[0] ;
 wire \sw_094_module_data_in[1] ;
 wire \sw_094_module_data_in[2] ;
 wire \sw_094_module_data_in[3] ;
 wire \sw_094_module_data_in[4] ;
 wire \sw_094_module_data_in[5] ;
 wire \sw_094_module_data_in[6] ;
 wire \sw_094_module_data_in[7] ;
 wire \sw_094_module_data_out[0] ;
 wire \sw_094_module_data_out[1] ;
 wire \sw_094_module_data_out[2] ;
 wire \sw_094_module_data_out[3] ;
 wire \sw_094_module_data_out[4] ;
 wire \sw_094_module_data_out[5] ;
 wire \sw_094_module_data_out[6] ;
 wire \sw_094_module_data_out[7] ;
 wire sw_094_scan_out;
 wire sw_095_clk_out;
 wire sw_095_data_out;
 wire sw_095_latch_out;
 wire \sw_095_module_data_in[0] ;
 wire \sw_095_module_data_in[1] ;
 wire \sw_095_module_data_in[2] ;
 wire \sw_095_module_data_in[3] ;
 wire \sw_095_module_data_in[4] ;
 wire \sw_095_module_data_in[5] ;
 wire \sw_095_module_data_in[6] ;
 wire \sw_095_module_data_in[7] ;
 wire \sw_095_module_data_out[0] ;
 wire \sw_095_module_data_out[1] ;
 wire \sw_095_module_data_out[2] ;
 wire \sw_095_module_data_out[3] ;
 wire \sw_095_module_data_out[4] ;
 wire \sw_095_module_data_out[5] ;
 wire \sw_095_module_data_out[6] ;
 wire \sw_095_module_data_out[7] ;
 wire sw_095_scan_out;
 wire sw_096_clk_out;
 wire sw_096_data_out;
 wire sw_096_latch_out;
 wire \sw_096_module_data_in[0] ;
 wire \sw_096_module_data_in[1] ;
 wire \sw_096_module_data_in[2] ;
 wire \sw_096_module_data_in[3] ;
 wire \sw_096_module_data_in[4] ;
 wire \sw_096_module_data_in[5] ;
 wire \sw_096_module_data_in[6] ;
 wire \sw_096_module_data_in[7] ;
 wire \sw_096_module_data_out[0] ;
 wire \sw_096_module_data_out[1] ;
 wire \sw_096_module_data_out[2] ;
 wire \sw_096_module_data_out[3] ;
 wire \sw_096_module_data_out[4] ;
 wire \sw_096_module_data_out[5] ;
 wire \sw_096_module_data_out[6] ;
 wire \sw_096_module_data_out[7] ;
 wire sw_096_scan_out;
 wire sw_097_clk_out;
 wire sw_097_data_out;
 wire sw_097_latch_out;
 wire \sw_097_module_data_in[0] ;
 wire \sw_097_module_data_in[1] ;
 wire \sw_097_module_data_in[2] ;
 wire \sw_097_module_data_in[3] ;
 wire \sw_097_module_data_in[4] ;
 wire \sw_097_module_data_in[5] ;
 wire \sw_097_module_data_in[6] ;
 wire \sw_097_module_data_in[7] ;
 wire \sw_097_module_data_out[0] ;
 wire \sw_097_module_data_out[1] ;
 wire \sw_097_module_data_out[2] ;
 wire \sw_097_module_data_out[3] ;
 wire \sw_097_module_data_out[4] ;
 wire \sw_097_module_data_out[5] ;
 wire \sw_097_module_data_out[6] ;
 wire \sw_097_module_data_out[7] ;
 wire sw_097_scan_out;
 wire sw_098_clk_out;
 wire sw_098_data_out;
 wire sw_098_latch_out;
 wire \sw_098_module_data_in[0] ;
 wire \sw_098_module_data_in[1] ;
 wire \sw_098_module_data_in[2] ;
 wire \sw_098_module_data_in[3] ;
 wire \sw_098_module_data_in[4] ;
 wire \sw_098_module_data_in[5] ;
 wire \sw_098_module_data_in[6] ;
 wire \sw_098_module_data_in[7] ;
 wire \sw_098_module_data_out[0] ;
 wire \sw_098_module_data_out[1] ;
 wire \sw_098_module_data_out[2] ;
 wire \sw_098_module_data_out[3] ;
 wire \sw_098_module_data_out[4] ;
 wire \sw_098_module_data_out[5] ;
 wire \sw_098_module_data_out[6] ;
 wire \sw_098_module_data_out[7] ;
 wire sw_098_scan_out;
 wire sw_099_clk_out;
 wire sw_099_data_out;
 wire sw_099_latch_out;
 wire \sw_099_module_data_in[0] ;
 wire \sw_099_module_data_in[1] ;
 wire \sw_099_module_data_in[2] ;
 wire \sw_099_module_data_in[3] ;
 wire \sw_099_module_data_in[4] ;
 wire \sw_099_module_data_in[5] ;
 wire \sw_099_module_data_in[6] ;
 wire \sw_099_module_data_in[7] ;
 wire \sw_099_module_data_out[0] ;
 wire \sw_099_module_data_out[1] ;
 wire \sw_099_module_data_out[2] ;
 wire \sw_099_module_data_out[3] ;
 wire \sw_099_module_data_out[4] ;
 wire \sw_099_module_data_out[5] ;
 wire \sw_099_module_data_out[6] ;
 wire \sw_099_module_data_out[7] ;
 wire sw_099_scan_out;
 wire sw_100_clk_out;
 wire sw_100_data_out;
 wire sw_100_latch_out;
 wire \sw_100_module_data_in[0] ;
 wire \sw_100_module_data_in[1] ;
 wire \sw_100_module_data_in[2] ;
 wire \sw_100_module_data_in[3] ;
 wire \sw_100_module_data_in[4] ;
 wire \sw_100_module_data_in[5] ;
 wire \sw_100_module_data_in[6] ;
 wire \sw_100_module_data_in[7] ;
 wire \sw_100_module_data_out[0] ;
 wire \sw_100_module_data_out[1] ;
 wire \sw_100_module_data_out[2] ;
 wire \sw_100_module_data_out[3] ;
 wire \sw_100_module_data_out[4] ;
 wire \sw_100_module_data_out[5] ;
 wire \sw_100_module_data_out[6] ;
 wire \sw_100_module_data_out[7] ;
 wire sw_100_scan_out;
 wire sw_101_clk_out;
 wire sw_101_data_out;
 wire sw_101_latch_out;
 wire \sw_101_module_data_in[0] ;
 wire \sw_101_module_data_in[1] ;
 wire \sw_101_module_data_in[2] ;
 wire \sw_101_module_data_in[3] ;
 wire \sw_101_module_data_in[4] ;
 wire \sw_101_module_data_in[5] ;
 wire \sw_101_module_data_in[6] ;
 wire \sw_101_module_data_in[7] ;
 wire \sw_101_module_data_out[0] ;
 wire \sw_101_module_data_out[1] ;
 wire \sw_101_module_data_out[2] ;
 wire \sw_101_module_data_out[3] ;
 wire \sw_101_module_data_out[4] ;
 wire \sw_101_module_data_out[5] ;
 wire \sw_101_module_data_out[6] ;
 wire \sw_101_module_data_out[7] ;
 wire sw_101_scan_out;
 wire sw_102_clk_out;
 wire sw_102_data_out;
 wire sw_102_latch_out;
 wire \sw_102_module_data_in[0] ;
 wire \sw_102_module_data_in[1] ;
 wire \sw_102_module_data_in[2] ;
 wire \sw_102_module_data_in[3] ;
 wire \sw_102_module_data_in[4] ;
 wire \sw_102_module_data_in[5] ;
 wire \sw_102_module_data_in[6] ;
 wire \sw_102_module_data_in[7] ;
 wire \sw_102_module_data_out[0] ;
 wire \sw_102_module_data_out[1] ;
 wire \sw_102_module_data_out[2] ;
 wire \sw_102_module_data_out[3] ;
 wire \sw_102_module_data_out[4] ;
 wire \sw_102_module_data_out[5] ;
 wire \sw_102_module_data_out[6] ;
 wire \sw_102_module_data_out[7] ;
 wire sw_102_scan_out;
 wire sw_103_clk_out;
 wire sw_103_data_out;
 wire sw_103_latch_out;
 wire \sw_103_module_data_in[0] ;
 wire \sw_103_module_data_in[1] ;
 wire \sw_103_module_data_in[2] ;
 wire \sw_103_module_data_in[3] ;
 wire \sw_103_module_data_in[4] ;
 wire \sw_103_module_data_in[5] ;
 wire \sw_103_module_data_in[6] ;
 wire \sw_103_module_data_in[7] ;
 wire \sw_103_module_data_out[0] ;
 wire \sw_103_module_data_out[1] ;
 wire \sw_103_module_data_out[2] ;
 wire \sw_103_module_data_out[3] ;
 wire \sw_103_module_data_out[4] ;
 wire \sw_103_module_data_out[5] ;
 wire \sw_103_module_data_out[6] ;
 wire \sw_103_module_data_out[7] ;
 wire sw_103_scan_out;
 wire sw_104_clk_out;
 wire sw_104_data_out;
 wire sw_104_latch_out;
 wire \sw_104_module_data_in[0] ;
 wire \sw_104_module_data_in[1] ;
 wire \sw_104_module_data_in[2] ;
 wire \sw_104_module_data_in[3] ;
 wire \sw_104_module_data_in[4] ;
 wire \sw_104_module_data_in[5] ;
 wire \sw_104_module_data_in[6] ;
 wire \sw_104_module_data_in[7] ;
 wire \sw_104_module_data_out[0] ;
 wire \sw_104_module_data_out[1] ;
 wire \sw_104_module_data_out[2] ;
 wire \sw_104_module_data_out[3] ;
 wire \sw_104_module_data_out[4] ;
 wire \sw_104_module_data_out[5] ;
 wire \sw_104_module_data_out[6] ;
 wire \sw_104_module_data_out[7] ;
 wire sw_104_scan_out;
 wire sw_105_clk_out;
 wire sw_105_data_out;
 wire sw_105_latch_out;
 wire \sw_105_module_data_in[0] ;
 wire \sw_105_module_data_in[1] ;
 wire \sw_105_module_data_in[2] ;
 wire \sw_105_module_data_in[3] ;
 wire \sw_105_module_data_in[4] ;
 wire \sw_105_module_data_in[5] ;
 wire \sw_105_module_data_in[6] ;
 wire \sw_105_module_data_in[7] ;
 wire \sw_105_module_data_out[0] ;
 wire \sw_105_module_data_out[1] ;
 wire \sw_105_module_data_out[2] ;
 wire \sw_105_module_data_out[3] ;
 wire \sw_105_module_data_out[4] ;
 wire \sw_105_module_data_out[5] ;
 wire \sw_105_module_data_out[6] ;
 wire \sw_105_module_data_out[7] ;
 wire sw_105_scan_out;
 wire sw_106_clk_out;
 wire sw_106_data_out;
 wire sw_106_latch_out;
 wire \sw_106_module_data_in[0] ;
 wire \sw_106_module_data_in[1] ;
 wire \sw_106_module_data_in[2] ;
 wire \sw_106_module_data_in[3] ;
 wire \sw_106_module_data_in[4] ;
 wire \sw_106_module_data_in[5] ;
 wire \sw_106_module_data_in[6] ;
 wire \sw_106_module_data_in[7] ;
 wire \sw_106_module_data_out[0] ;
 wire \sw_106_module_data_out[1] ;
 wire \sw_106_module_data_out[2] ;
 wire \sw_106_module_data_out[3] ;
 wire \sw_106_module_data_out[4] ;
 wire \sw_106_module_data_out[5] ;
 wire \sw_106_module_data_out[6] ;
 wire \sw_106_module_data_out[7] ;
 wire sw_106_scan_out;
 wire sw_107_clk_out;
 wire sw_107_data_out;
 wire sw_107_latch_out;
 wire \sw_107_module_data_in[0] ;
 wire \sw_107_module_data_in[1] ;
 wire \sw_107_module_data_in[2] ;
 wire \sw_107_module_data_in[3] ;
 wire \sw_107_module_data_in[4] ;
 wire \sw_107_module_data_in[5] ;
 wire \sw_107_module_data_in[6] ;
 wire \sw_107_module_data_in[7] ;
 wire \sw_107_module_data_out[0] ;
 wire \sw_107_module_data_out[1] ;
 wire \sw_107_module_data_out[2] ;
 wire \sw_107_module_data_out[3] ;
 wire \sw_107_module_data_out[4] ;
 wire \sw_107_module_data_out[5] ;
 wire \sw_107_module_data_out[6] ;
 wire \sw_107_module_data_out[7] ;
 wire sw_107_scan_out;
 wire sw_108_clk_out;
 wire sw_108_data_out;
 wire sw_108_latch_out;
 wire \sw_108_module_data_in[0] ;
 wire \sw_108_module_data_in[1] ;
 wire \sw_108_module_data_in[2] ;
 wire \sw_108_module_data_in[3] ;
 wire \sw_108_module_data_in[4] ;
 wire \sw_108_module_data_in[5] ;
 wire \sw_108_module_data_in[6] ;
 wire \sw_108_module_data_in[7] ;
 wire \sw_108_module_data_out[0] ;
 wire \sw_108_module_data_out[1] ;
 wire \sw_108_module_data_out[2] ;
 wire \sw_108_module_data_out[3] ;
 wire \sw_108_module_data_out[4] ;
 wire \sw_108_module_data_out[5] ;
 wire \sw_108_module_data_out[6] ;
 wire \sw_108_module_data_out[7] ;
 wire sw_108_scan_out;
 wire sw_109_clk_out;
 wire sw_109_data_out;
 wire sw_109_latch_out;
 wire \sw_109_module_data_in[0] ;
 wire \sw_109_module_data_in[1] ;
 wire \sw_109_module_data_in[2] ;
 wire \sw_109_module_data_in[3] ;
 wire \sw_109_module_data_in[4] ;
 wire \sw_109_module_data_in[5] ;
 wire \sw_109_module_data_in[6] ;
 wire \sw_109_module_data_in[7] ;
 wire \sw_109_module_data_out[0] ;
 wire \sw_109_module_data_out[1] ;
 wire \sw_109_module_data_out[2] ;
 wire \sw_109_module_data_out[3] ;
 wire \sw_109_module_data_out[4] ;
 wire \sw_109_module_data_out[5] ;
 wire \sw_109_module_data_out[6] ;
 wire \sw_109_module_data_out[7] ;
 wire sw_109_scan_out;
 wire sw_110_clk_out;
 wire sw_110_data_out;
 wire sw_110_latch_out;
 wire \sw_110_module_data_in[0] ;
 wire \sw_110_module_data_in[1] ;
 wire \sw_110_module_data_in[2] ;
 wire \sw_110_module_data_in[3] ;
 wire \sw_110_module_data_in[4] ;
 wire \sw_110_module_data_in[5] ;
 wire \sw_110_module_data_in[6] ;
 wire \sw_110_module_data_in[7] ;
 wire \sw_110_module_data_out[0] ;
 wire \sw_110_module_data_out[1] ;
 wire \sw_110_module_data_out[2] ;
 wire \sw_110_module_data_out[3] ;
 wire \sw_110_module_data_out[4] ;
 wire \sw_110_module_data_out[5] ;
 wire \sw_110_module_data_out[6] ;
 wire \sw_110_module_data_out[7] ;
 wire sw_110_scan_out;
 wire sw_111_clk_out;
 wire sw_111_data_out;
 wire sw_111_latch_out;
 wire \sw_111_module_data_in[0] ;
 wire \sw_111_module_data_in[1] ;
 wire \sw_111_module_data_in[2] ;
 wire \sw_111_module_data_in[3] ;
 wire \sw_111_module_data_in[4] ;
 wire \sw_111_module_data_in[5] ;
 wire \sw_111_module_data_in[6] ;
 wire \sw_111_module_data_in[7] ;
 wire \sw_111_module_data_out[0] ;
 wire \sw_111_module_data_out[1] ;
 wire \sw_111_module_data_out[2] ;
 wire \sw_111_module_data_out[3] ;
 wire \sw_111_module_data_out[4] ;
 wire \sw_111_module_data_out[5] ;
 wire \sw_111_module_data_out[6] ;
 wire \sw_111_module_data_out[7] ;
 wire sw_111_scan_out;
 wire sw_112_clk_out;
 wire sw_112_data_out;
 wire sw_112_latch_out;
 wire \sw_112_module_data_in[0] ;
 wire \sw_112_module_data_in[1] ;
 wire \sw_112_module_data_in[2] ;
 wire \sw_112_module_data_in[3] ;
 wire \sw_112_module_data_in[4] ;
 wire \sw_112_module_data_in[5] ;
 wire \sw_112_module_data_in[6] ;
 wire \sw_112_module_data_in[7] ;
 wire \sw_112_module_data_out[0] ;
 wire \sw_112_module_data_out[1] ;
 wire \sw_112_module_data_out[2] ;
 wire \sw_112_module_data_out[3] ;
 wire \sw_112_module_data_out[4] ;
 wire \sw_112_module_data_out[5] ;
 wire \sw_112_module_data_out[6] ;
 wire \sw_112_module_data_out[7] ;
 wire sw_112_scan_out;
 wire sw_113_clk_out;
 wire sw_113_data_out;
 wire sw_113_latch_out;
 wire \sw_113_module_data_in[0] ;
 wire \sw_113_module_data_in[1] ;
 wire \sw_113_module_data_in[2] ;
 wire \sw_113_module_data_in[3] ;
 wire \sw_113_module_data_in[4] ;
 wire \sw_113_module_data_in[5] ;
 wire \sw_113_module_data_in[6] ;
 wire \sw_113_module_data_in[7] ;
 wire \sw_113_module_data_out[0] ;
 wire \sw_113_module_data_out[1] ;
 wire \sw_113_module_data_out[2] ;
 wire \sw_113_module_data_out[3] ;
 wire \sw_113_module_data_out[4] ;
 wire \sw_113_module_data_out[5] ;
 wire \sw_113_module_data_out[6] ;
 wire \sw_113_module_data_out[7] ;
 wire sw_113_scan_out;
 wire sw_114_clk_out;
 wire sw_114_data_out;
 wire sw_114_latch_out;
 wire \sw_114_module_data_in[0] ;
 wire \sw_114_module_data_in[1] ;
 wire \sw_114_module_data_in[2] ;
 wire \sw_114_module_data_in[3] ;
 wire \sw_114_module_data_in[4] ;
 wire \sw_114_module_data_in[5] ;
 wire \sw_114_module_data_in[6] ;
 wire \sw_114_module_data_in[7] ;
 wire \sw_114_module_data_out[0] ;
 wire \sw_114_module_data_out[1] ;
 wire \sw_114_module_data_out[2] ;
 wire \sw_114_module_data_out[3] ;
 wire \sw_114_module_data_out[4] ;
 wire \sw_114_module_data_out[5] ;
 wire \sw_114_module_data_out[6] ;
 wire \sw_114_module_data_out[7] ;
 wire sw_114_scan_out;
 wire sw_115_clk_out;
 wire sw_115_data_out;
 wire sw_115_latch_out;
 wire \sw_115_module_data_in[0] ;
 wire \sw_115_module_data_in[1] ;
 wire \sw_115_module_data_in[2] ;
 wire \sw_115_module_data_in[3] ;
 wire \sw_115_module_data_in[4] ;
 wire \sw_115_module_data_in[5] ;
 wire \sw_115_module_data_in[6] ;
 wire \sw_115_module_data_in[7] ;
 wire \sw_115_module_data_out[0] ;
 wire \sw_115_module_data_out[1] ;
 wire \sw_115_module_data_out[2] ;
 wire \sw_115_module_data_out[3] ;
 wire \sw_115_module_data_out[4] ;
 wire \sw_115_module_data_out[5] ;
 wire \sw_115_module_data_out[6] ;
 wire \sw_115_module_data_out[7] ;
 wire sw_115_scan_out;
 wire sw_116_clk_out;
 wire sw_116_data_out;
 wire sw_116_latch_out;
 wire \sw_116_module_data_in[0] ;
 wire \sw_116_module_data_in[1] ;
 wire \sw_116_module_data_in[2] ;
 wire \sw_116_module_data_in[3] ;
 wire \sw_116_module_data_in[4] ;
 wire \sw_116_module_data_in[5] ;
 wire \sw_116_module_data_in[6] ;
 wire \sw_116_module_data_in[7] ;
 wire \sw_116_module_data_out[0] ;
 wire \sw_116_module_data_out[1] ;
 wire \sw_116_module_data_out[2] ;
 wire \sw_116_module_data_out[3] ;
 wire \sw_116_module_data_out[4] ;
 wire \sw_116_module_data_out[5] ;
 wire \sw_116_module_data_out[6] ;
 wire \sw_116_module_data_out[7] ;
 wire sw_116_scan_out;
 wire sw_117_clk_out;
 wire sw_117_data_out;
 wire sw_117_latch_out;
 wire \sw_117_module_data_in[0] ;
 wire \sw_117_module_data_in[1] ;
 wire \sw_117_module_data_in[2] ;
 wire \sw_117_module_data_in[3] ;
 wire \sw_117_module_data_in[4] ;
 wire \sw_117_module_data_in[5] ;
 wire \sw_117_module_data_in[6] ;
 wire \sw_117_module_data_in[7] ;
 wire \sw_117_module_data_out[0] ;
 wire \sw_117_module_data_out[1] ;
 wire \sw_117_module_data_out[2] ;
 wire \sw_117_module_data_out[3] ;
 wire \sw_117_module_data_out[4] ;
 wire \sw_117_module_data_out[5] ;
 wire \sw_117_module_data_out[6] ;
 wire \sw_117_module_data_out[7] ;
 wire sw_117_scan_out;
 wire sw_118_clk_out;
 wire sw_118_data_out;
 wire sw_118_latch_out;
 wire \sw_118_module_data_in[0] ;
 wire \sw_118_module_data_in[1] ;
 wire \sw_118_module_data_in[2] ;
 wire \sw_118_module_data_in[3] ;
 wire \sw_118_module_data_in[4] ;
 wire \sw_118_module_data_in[5] ;
 wire \sw_118_module_data_in[6] ;
 wire \sw_118_module_data_in[7] ;
 wire \sw_118_module_data_out[0] ;
 wire \sw_118_module_data_out[1] ;
 wire \sw_118_module_data_out[2] ;
 wire \sw_118_module_data_out[3] ;
 wire \sw_118_module_data_out[4] ;
 wire \sw_118_module_data_out[5] ;
 wire \sw_118_module_data_out[6] ;
 wire \sw_118_module_data_out[7] ;
 wire sw_118_scan_out;
 wire sw_119_clk_out;
 wire sw_119_data_out;
 wire sw_119_latch_out;
 wire \sw_119_module_data_in[0] ;
 wire \sw_119_module_data_in[1] ;
 wire \sw_119_module_data_in[2] ;
 wire \sw_119_module_data_in[3] ;
 wire \sw_119_module_data_in[4] ;
 wire \sw_119_module_data_in[5] ;
 wire \sw_119_module_data_in[6] ;
 wire \sw_119_module_data_in[7] ;
 wire \sw_119_module_data_out[0] ;
 wire \sw_119_module_data_out[1] ;
 wire \sw_119_module_data_out[2] ;
 wire \sw_119_module_data_out[3] ;
 wire \sw_119_module_data_out[4] ;
 wire \sw_119_module_data_out[5] ;
 wire \sw_119_module_data_out[6] ;
 wire \sw_119_module_data_out[7] ;
 wire sw_119_scan_out;
 wire sw_120_clk_out;
 wire sw_120_data_out;
 wire sw_120_latch_out;
 wire \sw_120_module_data_in[0] ;
 wire \sw_120_module_data_in[1] ;
 wire \sw_120_module_data_in[2] ;
 wire \sw_120_module_data_in[3] ;
 wire \sw_120_module_data_in[4] ;
 wire \sw_120_module_data_in[5] ;
 wire \sw_120_module_data_in[6] ;
 wire \sw_120_module_data_in[7] ;
 wire \sw_120_module_data_out[0] ;
 wire \sw_120_module_data_out[1] ;
 wire \sw_120_module_data_out[2] ;
 wire \sw_120_module_data_out[3] ;
 wire \sw_120_module_data_out[4] ;
 wire \sw_120_module_data_out[5] ;
 wire \sw_120_module_data_out[6] ;
 wire \sw_120_module_data_out[7] ;
 wire sw_120_scan_out;
 wire sw_121_clk_out;
 wire sw_121_data_out;
 wire sw_121_latch_out;
 wire \sw_121_module_data_in[0] ;
 wire \sw_121_module_data_in[1] ;
 wire \sw_121_module_data_in[2] ;
 wire \sw_121_module_data_in[3] ;
 wire \sw_121_module_data_in[4] ;
 wire \sw_121_module_data_in[5] ;
 wire \sw_121_module_data_in[6] ;
 wire \sw_121_module_data_in[7] ;
 wire \sw_121_module_data_out[0] ;
 wire \sw_121_module_data_out[1] ;
 wire \sw_121_module_data_out[2] ;
 wire \sw_121_module_data_out[3] ;
 wire \sw_121_module_data_out[4] ;
 wire \sw_121_module_data_out[5] ;
 wire \sw_121_module_data_out[6] ;
 wire \sw_121_module_data_out[7] ;
 wire sw_121_scan_out;
 wire sw_122_clk_out;
 wire sw_122_data_out;
 wire sw_122_latch_out;
 wire \sw_122_module_data_in[0] ;
 wire \sw_122_module_data_in[1] ;
 wire \sw_122_module_data_in[2] ;
 wire \sw_122_module_data_in[3] ;
 wire \sw_122_module_data_in[4] ;
 wire \sw_122_module_data_in[5] ;
 wire \sw_122_module_data_in[6] ;
 wire \sw_122_module_data_in[7] ;
 wire \sw_122_module_data_out[0] ;
 wire \sw_122_module_data_out[1] ;
 wire \sw_122_module_data_out[2] ;
 wire \sw_122_module_data_out[3] ;
 wire \sw_122_module_data_out[4] ;
 wire \sw_122_module_data_out[5] ;
 wire \sw_122_module_data_out[6] ;
 wire \sw_122_module_data_out[7] ;
 wire sw_122_scan_out;
 wire sw_123_clk_out;
 wire sw_123_data_out;
 wire sw_123_latch_out;
 wire \sw_123_module_data_in[0] ;
 wire \sw_123_module_data_in[1] ;
 wire \sw_123_module_data_in[2] ;
 wire \sw_123_module_data_in[3] ;
 wire \sw_123_module_data_in[4] ;
 wire \sw_123_module_data_in[5] ;
 wire \sw_123_module_data_in[6] ;
 wire \sw_123_module_data_in[7] ;
 wire \sw_123_module_data_out[0] ;
 wire \sw_123_module_data_out[1] ;
 wire \sw_123_module_data_out[2] ;
 wire \sw_123_module_data_out[3] ;
 wire \sw_123_module_data_out[4] ;
 wire \sw_123_module_data_out[5] ;
 wire \sw_123_module_data_out[6] ;
 wire \sw_123_module_data_out[7] ;
 wire sw_123_scan_out;
 wire sw_124_clk_out;
 wire sw_124_data_out;
 wire sw_124_latch_out;
 wire \sw_124_module_data_in[0] ;
 wire \sw_124_module_data_in[1] ;
 wire \sw_124_module_data_in[2] ;
 wire \sw_124_module_data_in[3] ;
 wire \sw_124_module_data_in[4] ;
 wire \sw_124_module_data_in[5] ;
 wire \sw_124_module_data_in[6] ;
 wire \sw_124_module_data_in[7] ;
 wire \sw_124_module_data_out[0] ;
 wire \sw_124_module_data_out[1] ;
 wire \sw_124_module_data_out[2] ;
 wire \sw_124_module_data_out[3] ;
 wire \sw_124_module_data_out[4] ;
 wire \sw_124_module_data_out[5] ;
 wire \sw_124_module_data_out[6] ;
 wire \sw_124_module_data_out[7] ;
 wire sw_124_scan_out;
 wire sw_125_clk_out;
 wire sw_125_data_out;
 wire sw_125_latch_out;
 wire \sw_125_module_data_in[0] ;
 wire \sw_125_module_data_in[1] ;
 wire \sw_125_module_data_in[2] ;
 wire \sw_125_module_data_in[3] ;
 wire \sw_125_module_data_in[4] ;
 wire \sw_125_module_data_in[5] ;
 wire \sw_125_module_data_in[6] ;
 wire \sw_125_module_data_in[7] ;
 wire \sw_125_module_data_out[0] ;
 wire \sw_125_module_data_out[1] ;
 wire \sw_125_module_data_out[2] ;
 wire \sw_125_module_data_out[3] ;
 wire \sw_125_module_data_out[4] ;
 wire \sw_125_module_data_out[5] ;
 wire \sw_125_module_data_out[6] ;
 wire \sw_125_module_data_out[7] ;
 wire sw_125_scan_out;
 wire sw_126_clk_out;
 wire sw_126_data_out;
 wire sw_126_latch_out;
 wire \sw_126_module_data_in[0] ;
 wire \sw_126_module_data_in[1] ;
 wire \sw_126_module_data_in[2] ;
 wire \sw_126_module_data_in[3] ;
 wire \sw_126_module_data_in[4] ;
 wire \sw_126_module_data_in[5] ;
 wire \sw_126_module_data_in[6] ;
 wire \sw_126_module_data_in[7] ;
 wire \sw_126_module_data_out[0] ;
 wire \sw_126_module_data_out[1] ;
 wire \sw_126_module_data_out[2] ;
 wire \sw_126_module_data_out[3] ;
 wire \sw_126_module_data_out[4] ;
 wire \sw_126_module_data_out[5] ;
 wire \sw_126_module_data_out[6] ;
 wire \sw_126_module_data_out[7] ;
 wire sw_126_scan_out;
 wire sw_127_clk_out;
 wire sw_127_data_out;
 wire sw_127_latch_out;
 wire \sw_127_module_data_in[0] ;
 wire \sw_127_module_data_in[1] ;
 wire \sw_127_module_data_in[2] ;
 wire \sw_127_module_data_in[3] ;
 wire \sw_127_module_data_in[4] ;
 wire \sw_127_module_data_in[5] ;
 wire \sw_127_module_data_in[6] ;
 wire \sw_127_module_data_in[7] ;
 wire \sw_127_module_data_out[0] ;
 wire \sw_127_module_data_out[1] ;
 wire \sw_127_module_data_out[2] ;
 wire \sw_127_module_data_out[3] ;
 wire \sw_127_module_data_out[4] ;
 wire \sw_127_module_data_out[5] ;
 wire \sw_127_module_data_out[6] ;
 wire \sw_127_module_data_out[7] ;
 wire sw_127_scan_out;
 wire sw_128_clk_out;
 wire sw_128_data_out;
 wire sw_128_latch_out;
 wire \sw_128_module_data_in[0] ;
 wire \sw_128_module_data_in[1] ;
 wire \sw_128_module_data_in[2] ;
 wire \sw_128_module_data_in[3] ;
 wire \sw_128_module_data_in[4] ;
 wire \sw_128_module_data_in[5] ;
 wire \sw_128_module_data_in[6] ;
 wire \sw_128_module_data_in[7] ;
 wire \sw_128_module_data_out[0] ;
 wire \sw_128_module_data_out[1] ;
 wire \sw_128_module_data_out[2] ;
 wire \sw_128_module_data_out[3] ;
 wire \sw_128_module_data_out[4] ;
 wire \sw_128_module_data_out[5] ;
 wire \sw_128_module_data_out[6] ;
 wire \sw_128_module_data_out[7] ;
 wire sw_128_scan_out;
 wire sw_129_clk_out;
 wire sw_129_data_out;
 wire sw_129_latch_out;
 wire \sw_129_module_data_in[0] ;
 wire \sw_129_module_data_in[1] ;
 wire \sw_129_module_data_in[2] ;
 wire \sw_129_module_data_in[3] ;
 wire \sw_129_module_data_in[4] ;
 wire \sw_129_module_data_in[5] ;
 wire \sw_129_module_data_in[6] ;
 wire \sw_129_module_data_in[7] ;
 wire \sw_129_module_data_out[0] ;
 wire \sw_129_module_data_out[1] ;
 wire \sw_129_module_data_out[2] ;
 wire \sw_129_module_data_out[3] ;
 wire \sw_129_module_data_out[4] ;
 wire \sw_129_module_data_out[5] ;
 wire \sw_129_module_data_out[6] ;
 wire \sw_129_module_data_out[7] ;
 wire sw_129_scan_out;
 wire sw_130_clk_out;
 wire sw_130_data_out;
 wire sw_130_latch_out;
 wire \sw_130_module_data_in[0] ;
 wire \sw_130_module_data_in[1] ;
 wire \sw_130_module_data_in[2] ;
 wire \sw_130_module_data_in[3] ;
 wire \sw_130_module_data_in[4] ;
 wire \sw_130_module_data_in[5] ;
 wire \sw_130_module_data_in[6] ;
 wire \sw_130_module_data_in[7] ;
 wire \sw_130_module_data_out[0] ;
 wire \sw_130_module_data_out[1] ;
 wire \sw_130_module_data_out[2] ;
 wire \sw_130_module_data_out[3] ;
 wire \sw_130_module_data_out[4] ;
 wire \sw_130_module_data_out[5] ;
 wire \sw_130_module_data_out[6] ;
 wire \sw_130_module_data_out[7] ;
 wire sw_130_scan_out;
 wire sw_131_clk_out;
 wire sw_131_data_out;
 wire sw_131_latch_out;
 wire \sw_131_module_data_in[0] ;
 wire \sw_131_module_data_in[1] ;
 wire \sw_131_module_data_in[2] ;
 wire \sw_131_module_data_in[3] ;
 wire \sw_131_module_data_in[4] ;
 wire \sw_131_module_data_in[5] ;
 wire \sw_131_module_data_in[6] ;
 wire \sw_131_module_data_in[7] ;
 wire \sw_131_module_data_out[0] ;
 wire \sw_131_module_data_out[1] ;
 wire \sw_131_module_data_out[2] ;
 wire \sw_131_module_data_out[3] ;
 wire \sw_131_module_data_out[4] ;
 wire \sw_131_module_data_out[5] ;
 wire \sw_131_module_data_out[6] ;
 wire \sw_131_module_data_out[7] ;
 wire sw_131_scan_out;
 wire sw_132_clk_out;
 wire sw_132_data_out;
 wire sw_132_latch_out;
 wire \sw_132_module_data_in[0] ;
 wire \sw_132_module_data_in[1] ;
 wire \sw_132_module_data_in[2] ;
 wire \sw_132_module_data_in[3] ;
 wire \sw_132_module_data_in[4] ;
 wire \sw_132_module_data_in[5] ;
 wire \sw_132_module_data_in[6] ;
 wire \sw_132_module_data_in[7] ;
 wire \sw_132_module_data_out[0] ;
 wire \sw_132_module_data_out[1] ;
 wire \sw_132_module_data_out[2] ;
 wire \sw_132_module_data_out[3] ;
 wire \sw_132_module_data_out[4] ;
 wire \sw_132_module_data_out[5] ;
 wire \sw_132_module_data_out[6] ;
 wire \sw_132_module_data_out[7] ;
 wire sw_132_scan_out;
 wire sw_133_clk_out;
 wire sw_133_data_out;
 wire sw_133_latch_out;
 wire \sw_133_module_data_in[0] ;
 wire \sw_133_module_data_in[1] ;
 wire \sw_133_module_data_in[2] ;
 wire \sw_133_module_data_in[3] ;
 wire \sw_133_module_data_in[4] ;
 wire \sw_133_module_data_in[5] ;
 wire \sw_133_module_data_in[6] ;
 wire \sw_133_module_data_in[7] ;
 wire \sw_133_module_data_out[0] ;
 wire \sw_133_module_data_out[1] ;
 wire \sw_133_module_data_out[2] ;
 wire \sw_133_module_data_out[3] ;
 wire \sw_133_module_data_out[4] ;
 wire \sw_133_module_data_out[5] ;
 wire \sw_133_module_data_out[6] ;
 wire \sw_133_module_data_out[7] ;
 wire sw_133_scan_out;
 wire sw_134_clk_out;
 wire sw_134_data_out;
 wire sw_134_latch_out;
 wire \sw_134_module_data_in[0] ;
 wire \sw_134_module_data_in[1] ;
 wire \sw_134_module_data_in[2] ;
 wire \sw_134_module_data_in[3] ;
 wire \sw_134_module_data_in[4] ;
 wire \sw_134_module_data_in[5] ;
 wire \sw_134_module_data_in[6] ;
 wire \sw_134_module_data_in[7] ;
 wire \sw_134_module_data_out[0] ;
 wire \sw_134_module_data_out[1] ;
 wire \sw_134_module_data_out[2] ;
 wire \sw_134_module_data_out[3] ;
 wire \sw_134_module_data_out[4] ;
 wire \sw_134_module_data_out[5] ;
 wire \sw_134_module_data_out[6] ;
 wire \sw_134_module_data_out[7] ;
 wire sw_134_scan_out;
 wire sw_135_clk_out;
 wire sw_135_data_out;
 wire sw_135_latch_out;
 wire \sw_135_module_data_in[0] ;
 wire \sw_135_module_data_in[1] ;
 wire \sw_135_module_data_in[2] ;
 wire \sw_135_module_data_in[3] ;
 wire \sw_135_module_data_in[4] ;
 wire \sw_135_module_data_in[5] ;
 wire \sw_135_module_data_in[6] ;
 wire \sw_135_module_data_in[7] ;
 wire \sw_135_module_data_out[0] ;
 wire \sw_135_module_data_out[1] ;
 wire \sw_135_module_data_out[2] ;
 wire \sw_135_module_data_out[3] ;
 wire \sw_135_module_data_out[4] ;
 wire \sw_135_module_data_out[5] ;
 wire \sw_135_module_data_out[6] ;
 wire \sw_135_module_data_out[7] ;
 wire sw_135_scan_out;
 wire sw_136_clk_out;
 wire sw_136_data_out;
 wire sw_136_latch_out;
 wire \sw_136_module_data_in[0] ;
 wire \sw_136_module_data_in[1] ;
 wire \sw_136_module_data_in[2] ;
 wire \sw_136_module_data_in[3] ;
 wire \sw_136_module_data_in[4] ;
 wire \sw_136_module_data_in[5] ;
 wire \sw_136_module_data_in[6] ;
 wire \sw_136_module_data_in[7] ;
 wire \sw_136_module_data_out[0] ;
 wire \sw_136_module_data_out[1] ;
 wire \sw_136_module_data_out[2] ;
 wire \sw_136_module_data_out[3] ;
 wire \sw_136_module_data_out[4] ;
 wire \sw_136_module_data_out[5] ;
 wire \sw_136_module_data_out[6] ;
 wire \sw_136_module_data_out[7] ;
 wire sw_136_scan_out;
 wire sw_137_clk_out;
 wire sw_137_data_out;
 wire sw_137_latch_out;
 wire \sw_137_module_data_in[0] ;
 wire \sw_137_module_data_in[1] ;
 wire \sw_137_module_data_in[2] ;
 wire \sw_137_module_data_in[3] ;
 wire \sw_137_module_data_in[4] ;
 wire \sw_137_module_data_in[5] ;
 wire \sw_137_module_data_in[6] ;
 wire \sw_137_module_data_in[7] ;
 wire \sw_137_module_data_out[0] ;
 wire \sw_137_module_data_out[1] ;
 wire \sw_137_module_data_out[2] ;
 wire \sw_137_module_data_out[3] ;
 wire \sw_137_module_data_out[4] ;
 wire \sw_137_module_data_out[5] ;
 wire \sw_137_module_data_out[6] ;
 wire \sw_137_module_data_out[7] ;
 wire sw_137_scan_out;
 wire sw_138_clk_out;
 wire sw_138_data_out;
 wire sw_138_latch_out;
 wire \sw_138_module_data_in[0] ;
 wire \sw_138_module_data_in[1] ;
 wire \sw_138_module_data_in[2] ;
 wire \sw_138_module_data_in[3] ;
 wire \sw_138_module_data_in[4] ;
 wire \sw_138_module_data_in[5] ;
 wire \sw_138_module_data_in[6] ;
 wire \sw_138_module_data_in[7] ;
 wire \sw_138_module_data_out[0] ;
 wire \sw_138_module_data_out[1] ;
 wire \sw_138_module_data_out[2] ;
 wire \sw_138_module_data_out[3] ;
 wire \sw_138_module_data_out[4] ;
 wire \sw_138_module_data_out[5] ;
 wire \sw_138_module_data_out[6] ;
 wire \sw_138_module_data_out[7] ;
 wire sw_138_scan_out;
 wire sw_139_clk_out;
 wire sw_139_data_out;
 wire sw_139_latch_out;
 wire \sw_139_module_data_in[0] ;
 wire \sw_139_module_data_in[1] ;
 wire \sw_139_module_data_in[2] ;
 wire \sw_139_module_data_in[3] ;
 wire \sw_139_module_data_in[4] ;
 wire \sw_139_module_data_in[5] ;
 wire \sw_139_module_data_in[6] ;
 wire \sw_139_module_data_in[7] ;
 wire \sw_139_module_data_out[0] ;
 wire \sw_139_module_data_out[1] ;
 wire \sw_139_module_data_out[2] ;
 wire \sw_139_module_data_out[3] ;
 wire \sw_139_module_data_out[4] ;
 wire \sw_139_module_data_out[5] ;
 wire \sw_139_module_data_out[6] ;
 wire \sw_139_module_data_out[7] ;
 wire sw_139_scan_out;
 wire sw_140_clk_out;
 wire sw_140_data_out;
 wire sw_140_latch_out;
 wire \sw_140_module_data_in[0] ;
 wire \sw_140_module_data_in[1] ;
 wire \sw_140_module_data_in[2] ;
 wire \sw_140_module_data_in[3] ;
 wire \sw_140_module_data_in[4] ;
 wire \sw_140_module_data_in[5] ;
 wire \sw_140_module_data_in[6] ;
 wire \sw_140_module_data_in[7] ;
 wire \sw_140_module_data_out[0] ;
 wire \sw_140_module_data_out[1] ;
 wire \sw_140_module_data_out[2] ;
 wire \sw_140_module_data_out[3] ;
 wire \sw_140_module_data_out[4] ;
 wire \sw_140_module_data_out[5] ;
 wire \sw_140_module_data_out[6] ;
 wire \sw_140_module_data_out[7] ;
 wire sw_140_scan_out;
 wire sw_141_clk_out;
 wire sw_141_data_out;
 wire sw_141_latch_out;
 wire \sw_141_module_data_in[0] ;
 wire \sw_141_module_data_in[1] ;
 wire \sw_141_module_data_in[2] ;
 wire \sw_141_module_data_in[3] ;
 wire \sw_141_module_data_in[4] ;
 wire \sw_141_module_data_in[5] ;
 wire \sw_141_module_data_in[6] ;
 wire \sw_141_module_data_in[7] ;
 wire \sw_141_module_data_out[0] ;
 wire \sw_141_module_data_out[1] ;
 wire \sw_141_module_data_out[2] ;
 wire \sw_141_module_data_out[3] ;
 wire \sw_141_module_data_out[4] ;
 wire \sw_141_module_data_out[5] ;
 wire \sw_141_module_data_out[6] ;
 wire \sw_141_module_data_out[7] ;
 wire sw_141_scan_out;
 wire sw_142_clk_out;
 wire sw_142_data_out;
 wire sw_142_latch_out;
 wire \sw_142_module_data_in[0] ;
 wire \sw_142_module_data_in[1] ;
 wire \sw_142_module_data_in[2] ;
 wire \sw_142_module_data_in[3] ;
 wire \sw_142_module_data_in[4] ;
 wire \sw_142_module_data_in[5] ;
 wire \sw_142_module_data_in[6] ;
 wire \sw_142_module_data_in[7] ;
 wire \sw_142_module_data_out[0] ;
 wire \sw_142_module_data_out[1] ;
 wire \sw_142_module_data_out[2] ;
 wire \sw_142_module_data_out[3] ;
 wire \sw_142_module_data_out[4] ;
 wire \sw_142_module_data_out[5] ;
 wire \sw_142_module_data_out[6] ;
 wire \sw_142_module_data_out[7] ;
 wire sw_142_scan_out;
 wire sw_143_clk_out;
 wire sw_143_data_out;
 wire sw_143_latch_out;
 wire \sw_143_module_data_in[0] ;
 wire \sw_143_module_data_in[1] ;
 wire \sw_143_module_data_in[2] ;
 wire \sw_143_module_data_in[3] ;
 wire \sw_143_module_data_in[4] ;
 wire \sw_143_module_data_in[5] ;
 wire \sw_143_module_data_in[6] ;
 wire \sw_143_module_data_in[7] ;
 wire \sw_143_module_data_out[0] ;
 wire \sw_143_module_data_out[1] ;
 wire \sw_143_module_data_out[2] ;
 wire \sw_143_module_data_out[3] ;
 wire \sw_143_module_data_out[4] ;
 wire \sw_143_module_data_out[5] ;
 wire \sw_143_module_data_out[6] ;
 wire \sw_143_module_data_out[7] ;
 wire sw_143_scan_out;
 wire sw_144_clk_out;
 wire sw_144_data_out;
 wire sw_144_latch_out;
 wire \sw_144_module_data_in[0] ;
 wire \sw_144_module_data_in[1] ;
 wire \sw_144_module_data_in[2] ;
 wire \sw_144_module_data_in[3] ;
 wire \sw_144_module_data_in[4] ;
 wire \sw_144_module_data_in[5] ;
 wire \sw_144_module_data_in[6] ;
 wire \sw_144_module_data_in[7] ;
 wire \sw_144_module_data_out[0] ;
 wire \sw_144_module_data_out[1] ;
 wire \sw_144_module_data_out[2] ;
 wire \sw_144_module_data_out[3] ;
 wire \sw_144_module_data_out[4] ;
 wire \sw_144_module_data_out[5] ;
 wire \sw_144_module_data_out[6] ;
 wire \sw_144_module_data_out[7] ;
 wire sw_144_scan_out;
 wire sw_145_clk_out;
 wire sw_145_data_out;
 wire sw_145_latch_out;
 wire \sw_145_module_data_in[0] ;
 wire \sw_145_module_data_in[1] ;
 wire \sw_145_module_data_in[2] ;
 wire \sw_145_module_data_in[3] ;
 wire \sw_145_module_data_in[4] ;
 wire \sw_145_module_data_in[5] ;
 wire \sw_145_module_data_in[6] ;
 wire \sw_145_module_data_in[7] ;
 wire \sw_145_module_data_out[0] ;
 wire \sw_145_module_data_out[1] ;
 wire \sw_145_module_data_out[2] ;
 wire \sw_145_module_data_out[3] ;
 wire \sw_145_module_data_out[4] ;
 wire \sw_145_module_data_out[5] ;
 wire \sw_145_module_data_out[6] ;
 wire \sw_145_module_data_out[7] ;
 wire sw_145_scan_out;
 wire sw_146_clk_out;
 wire sw_146_data_out;
 wire sw_146_latch_out;
 wire \sw_146_module_data_in[0] ;
 wire \sw_146_module_data_in[1] ;
 wire \sw_146_module_data_in[2] ;
 wire \sw_146_module_data_in[3] ;
 wire \sw_146_module_data_in[4] ;
 wire \sw_146_module_data_in[5] ;
 wire \sw_146_module_data_in[6] ;
 wire \sw_146_module_data_in[7] ;
 wire \sw_146_module_data_out[0] ;
 wire \sw_146_module_data_out[1] ;
 wire \sw_146_module_data_out[2] ;
 wire \sw_146_module_data_out[3] ;
 wire \sw_146_module_data_out[4] ;
 wire \sw_146_module_data_out[5] ;
 wire \sw_146_module_data_out[6] ;
 wire \sw_146_module_data_out[7] ;
 wire sw_146_scan_out;
 wire sw_147_clk_out;
 wire sw_147_data_out;
 wire sw_147_latch_out;
 wire \sw_147_module_data_in[0] ;
 wire \sw_147_module_data_in[1] ;
 wire \sw_147_module_data_in[2] ;
 wire \sw_147_module_data_in[3] ;
 wire \sw_147_module_data_in[4] ;
 wire \sw_147_module_data_in[5] ;
 wire \sw_147_module_data_in[6] ;
 wire \sw_147_module_data_in[7] ;
 wire \sw_147_module_data_out[0] ;
 wire \sw_147_module_data_out[1] ;
 wire \sw_147_module_data_out[2] ;
 wire \sw_147_module_data_out[3] ;
 wire \sw_147_module_data_out[4] ;
 wire \sw_147_module_data_out[5] ;
 wire \sw_147_module_data_out[6] ;
 wire \sw_147_module_data_out[7] ;
 wire sw_147_scan_out;
 wire sw_148_clk_out;
 wire sw_148_data_out;
 wire sw_148_latch_out;
 wire \sw_148_module_data_in[0] ;
 wire \sw_148_module_data_in[1] ;
 wire \sw_148_module_data_in[2] ;
 wire \sw_148_module_data_in[3] ;
 wire \sw_148_module_data_in[4] ;
 wire \sw_148_module_data_in[5] ;
 wire \sw_148_module_data_in[6] ;
 wire \sw_148_module_data_in[7] ;
 wire \sw_148_module_data_out[0] ;
 wire \sw_148_module_data_out[1] ;
 wire \sw_148_module_data_out[2] ;
 wire \sw_148_module_data_out[3] ;
 wire \sw_148_module_data_out[4] ;
 wire \sw_148_module_data_out[5] ;
 wire \sw_148_module_data_out[6] ;
 wire \sw_148_module_data_out[7] ;
 wire sw_148_scan_out;
 wire sw_149_clk_out;
 wire sw_149_data_out;
 wire sw_149_latch_out;
 wire \sw_149_module_data_in[0] ;
 wire \sw_149_module_data_in[1] ;
 wire \sw_149_module_data_in[2] ;
 wire \sw_149_module_data_in[3] ;
 wire \sw_149_module_data_in[4] ;
 wire \sw_149_module_data_in[5] ;
 wire \sw_149_module_data_in[6] ;
 wire \sw_149_module_data_in[7] ;
 wire \sw_149_module_data_out[0] ;
 wire \sw_149_module_data_out[1] ;
 wire \sw_149_module_data_out[2] ;
 wire \sw_149_module_data_out[3] ;
 wire \sw_149_module_data_out[4] ;
 wire \sw_149_module_data_out[5] ;
 wire \sw_149_module_data_out[6] ;
 wire \sw_149_module_data_out[7] ;
 wire sw_149_scan_out;
 wire sw_150_clk_out;
 wire sw_150_data_out;
 wire sw_150_latch_out;
 wire \sw_150_module_data_in[0] ;
 wire \sw_150_module_data_in[1] ;
 wire \sw_150_module_data_in[2] ;
 wire \sw_150_module_data_in[3] ;
 wire \sw_150_module_data_in[4] ;
 wire \sw_150_module_data_in[5] ;
 wire \sw_150_module_data_in[6] ;
 wire \sw_150_module_data_in[7] ;
 wire \sw_150_module_data_out[0] ;
 wire \sw_150_module_data_out[1] ;
 wire \sw_150_module_data_out[2] ;
 wire \sw_150_module_data_out[3] ;
 wire \sw_150_module_data_out[4] ;
 wire \sw_150_module_data_out[5] ;
 wire \sw_150_module_data_out[6] ;
 wire \sw_150_module_data_out[7] ;
 wire sw_150_scan_out;
 wire sw_151_clk_out;
 wire sw_151_data_out;
 wire sw_151_latch_out;
 wire \sw_151_module_data_in[0] ;
 wire \sw_151_module_data_in[1] ;
 wire \sw_151_module_data_in[2] ;
 wire \sw_151_module_data_in[3] ;
 wire \sw_151_module_data_in[4] ;
 wire \sw_151_module_data_in[5] ;
 wire \sw_151_module_data_in[6] ;
 wire \sw_151_module_data_in[7] ;
 wire \sw_151_module_data_out[0] ;
 wire \sw_151_module_data_out[1] ;
 wire \sw_151_module_data_out[2] ;
 wire \sw_151_module_data_out[3] ;
 wire \sw_151_module_data_out[4] ;
 wire \sw_151_module_data_out[5] ;
 wire \sw_151_module_data_out[6] ;
 wire \sw_151_module_data_out[7] ;
 wire sw_151_scan_out;
 wire sw_152_clk_out;
 wire sw_152_data_out;
 wire sw_152_latch_out;
 wire \sw_152_module_data_in[0] ;
 wire \sw_152_module_data_in[1] ;
 wire \sw_152_module_data_in[2] ;
 wire \sw_152_module_data_in[3] ;
 wire \sw_152_module_data_in[4] ;
 wire \sw_152_module_data_in[5] ;
 wire \sw_152_module_data_in[6] ;
 wire \sw_152_module_data_in[7] ;
 wire \sw_152_module_data_out[0] ;
 wire \sw_152_module_data_out[1] ;
 wire \sw_152_module_data_out[2] ;
 wire \sw_152_module_data_out[3] ;
 wire \sw_152_module_data_out[4] ;
 wire \sw_152_module_data_out[5] ;
 wire \sw_152_module_data_out[6] ;
 wire \sw_152_module_data_out[7] ;
 wire sw_152_scan_out;
 wire sw_153_clk_out;
 wire sw_153_data_out;
 wire sw_153_latch_out;
 wire \sw_153_module_data_in[0] ;
 wire \sw_153_module_data_in[1] ;
 wire \sw_153_module_data_in[2] ;
 wire \sw_153_module_data_in[3] ;
 wire \sw_153_module_data_in[4] ;
 wire \sw_153_module_data_in[5] ;
 wire \sw_153_module_data_in[6] ;
 wire \sw_153_module_data_in[7] ;
 wire \sw_153_module_data_out[0] ;
 wire \sw_153_module_data_out[1] ;
 wire \sw_153_module_data_out[2] ;
 wire \sw_153_module_data_out[3] ;
 wire \sw_153_module_data_out[4] ;
 wire \sw_153_module_data_out[5] ;
 wire \sw_153_module_data_out[6] ;
 wire \sw_153_module_data_out[7] ;
 wire sw_153_scan_out;
 wire sw_154_clk_out;
 wire sw_154_data_out;
 wire sw_154_latch_out;
 wire \sw_154_module_data_in[0] ;
 wire \sw_154_module_data_in[1] ;
 wire \sw_154_module_data_in[2] ;
 wire \sw_154_module_data_in[3] ;
 wire \sw_154_module_data_in[4] ;
 wire \sw_154_module_data_in[5] ;
 wire \sw_154_module_data_in[6] ;
 wire \sw_154_module_data_in[7] ;
 wire \sw_154_module_data_out[0] ;
 wire \sw_154_module_data_out[1] ;
 wire \sw_154_module_data_out[2] ;
 wire \sw_154_module_data_out[3] ;
 wire \sw_154_module_data_out[4] ;
 wire \sw_154_module_data_out[5] ;
 wire \sw_154_module_data_out[6] ;
 wire \sw_154_module_data_out[7] ;
 wire sw_154_scan_out;
 wire sw_155_clk_out;
 wire sw_155_data_out;
 wire sw_155_latch_out;
 wire \sw_155_module_data_in[0] ;
 wire \sw_155_module_data_in[1] ;
 wire \sw_155_module_data_in[2] ;
 wire \sw_155_module_data_in[3] ;
 wire \sw_155_module_data_in[4] ;
 wire \sw_155_module_data_in[5] ;
 wire \sw_155_module_data_in[6] ;
 wire \sw_155_module_data_in[7] ;
 wire \sw_155_module_data_out[0] ;
 wire \sw_155_module_data_out[1] ;
 wire \sw_155_module_data_out[2] ;
 wire \sw_155_module_data_out[3] ;
 wire \sw_155_module_data_out[4] ;
 wire \sw_155_module_data_out[5] ;
 wire \sw_155_module_data_out[6] ;
 wire \sw_155_module_data_out[7] ;
 wire sw_155_scan_out;
 wire sw_156_clk_out;
 wire sw_156_data_out;
 wire sw_156_latch_out;
 wire \sw_156_module_data_in[0] ;
 wire \sw_156_module_data_in[1] ;
 wire \sw_156_module_data_in[2] ;
 wire \sw_156_module_data_in[3] ;
 wire \sw_156_module_data_in[4] ;
 wire \sw_156_module_data_in[5] ;
 wire \sw_156_module_data_in[6] ;
 wire \sw_156_module_data_in[7] ;
 wire \sw_156_module_data_out[0] ;
 wire \sw_156_module_data_out[1] ;
 wire \sw_156_module_data_out[2] ;
 wire \sw_156_module_data_out[3] ;
 wire \sw_156_module_data_out[4] ;
 wire \sw_156_module_data_out[5] ;
 wire \sw_156_module_data_out[6] ;
 wire \sw_156_module_data_out[7] ;
 wire sw_156_scan_out;
 wire sw_157_clk_out;
 wire sw_157_data_out;
 wire sw_157_latch_out;
 wire \sw_157_module_data_in[0] ;
 wire \sw_157_module_data_in[1] ;
 wire \sw_157_module_data_in[2] ;
 wire \sw_157_module_data_in[3] ;
 wire \sw_157_module_data_in[4] ;
 wire \sw_157_module_data_in[5] ;
 wire \sw_157_module_data_in[6] ;
 wire \sw_157_module_data_in[7] ;
 wire \sw_157_module_data_out[0] ;
 wire \sw_157_module_data_out[1] ;
 wire \sw_157_module_data_out[2] ;
 wire \sw_157_module_data_out[3] ;
 wire \sw_157_module_data_out[4] ;
 wire \sw_157_module_data_out[5] ;
 wire \sw_157_module_data_out[6] ;
 wire \sw_157_module_data_out[7] ;
 wire sw_157_scan_out;
 wire sw_158_clk_out;
 wire sw_158_data_out;
 wire sw_158_latch_out;
 wire \sw_158_module_data_in[0] ;
 wire \sw_158_module_data_in[1] ;
 wire \sw_158_module_data_in[2] ;
 wire \sw_158_module_data_in[3] ;
 wire \sw_158_module_data_in[4] ;
 wire \sw_158_module_data_in[5] ;
 wire \sw_158_module_data_in[6] ;
 wire \sw_158_module_data_in[7] ;
 wire \sw_158_module_data_out[0] ;
 wire \sw_158_module_data_out[1] ;
 wire \sw_158_module_data_out[2] ;
 wire \sw_158_module_data_out[3] ;
 wire \sw_158_module_data_out[4] ;
 wire \sw_158_module_data_out[5] ;
 wire \sw_158_module_data_out[6] ;
 wire \sw_158_module_data_out[7] ;
 wire sw_158_scan_out;
 wire sw_159_clk_out;
 wire sw_159_data_out;
 wire sw_159_latch_out;
 wire \sw_159_module_data_in[0] ;
 wire \sw_159_module_data_in[1] ;
 wire \sw_159_module_data_in[2] ;
 wire \sw_159_module_data_in[3] ;
 wire \sw_159_module_data_in[4] ;
 wire \sw_159_module_data_in[5] ;
 wire \sw_159_module_data_in[6] ;
 wire \sw_159_module_data_in[7] ;
 wire \sw_159_module_data_out[0] ;
 wire \sw_159_module_data_out[1] ;
 wire \sw_159_module_data_out[2] ;
 wire \sw_159_module_data_out[3] ;
 wire \sw_159_module_data_out[4] ;
 wire \sw_159_module_data_out[5] ;
 wire \sw_159_module_data_out[6] ;
 wire \sw_159_module_data_out[7] ;
 wire sw_159_scan_out;
 wire sw_160_clk_out;
 wire sw_160_data_out;
 wire sw_160_latch_out;
 wire \sw_160_module_data_in[0] ;
 wire \sw_160_module_data_in[1] ;
 wire \sw_160_module_data_in[2] ;
 wire \sw_160_module_data_in[3] ;
 wire \sw_160_module_data_in[4] ;
 wire \sw_160_module_data_in[5] ;
 wire \sw_160_module_data_in[6] ;
 wire \sw_160_module_data_in[7] ;
 wire \sw_160_module_data_out[0] ;
 wire \sw_160_module_data_out[1] ;
 wire \sw_160_module_data_out[2] ;
 wire \sw_160_module_data_out[3] ;
 wire \sw_160_module_data_out[4] ;
 wire \sw_160_module_data_out[5] ;
 wire \sw_160_module_data_out[6] ;
 wire \sw_160_module_data_out[7] ;
 wire sw_160_scan_out;
 wire sw_161_clk_out;
 wire sw_161_data_out;
 wire sw_161_latch_out;
 wire \sw_161_module_data_in[0] ;
 wire \sw_161_module_data_in[1] ;
 wire \sw_161_module_data_in[2] ;
 wire \sw_161_module_data_in[3] ;
 wire \sw_161_module_data_in[4] ;
 wire \sw_161_module_data_in[5] ;
 wire \sw_161_module_data_in[6] ;
 wire \sw_161_module_data_in[7] ;
 wire \sw_161_module_data_out[0] ;
 wire \sw_161_module_data_out[1] ;
 wire \sw_161_module_data_out[2] ;
 wire \sw_161_module_data_out[3] ;
 wire \sw_161_module_data_out[4] ;
 wire \sw_161_module_data_out[5] ;
 wire \sw_161_module_data_out[6] ;
 wire \sw_161_module_data_out[7] ;
 wire sw_161_scan_out;
 wire sw_162_clk_out;
 wire sw_162_data_out;
 wire sw_162_latch_out;
 wire \sw_162_module_data_in[0] ;
 wire \sw_162_module_data_in[1] ;
 wire \sw_162_module_data_in[2] ;
 wire \sw_162_module_data_in[3] ;
 wire \sw_162_module_data_in[4] ;
 wire \sw_162_module_data_in[5] ;
 wire \sw_162_module_data_in[6] ;
 wire \sw_162_module_data_in[7] ;
 wire \sw_162_module_data_out[0] ;
 wire \sw_162_module_data_out[1] ;
 wire \sw_162_module_data_out[2] ;
 wire \sw_162_module_data_out[3] ;
 wire \sw_162_module_data_out[4] ;
 wire \sw_162_module_data_out[5] ;
 wire \sw_162_module_data_out[6] ;
 wire \sw_162_module_data_out[7] ;
 wire sw_162_scan_out;
 wire sw_163_clk_out;
 wire sw_163_data_out;
 wire sw_163_latch_out;
 wire \sw_163_module_data_in[0] ;
 wire \sw_163_module_data_in[1] ;
 wire \sw_163_module_data_in[2] ;
 wire \sw_163_module_data_in[3] ;
 wire \sw_163_module_data_in[4] ;
 wire \sw_163_module_data_in[5] ;
 wire \sw_163_module_data_in[6] ;
 wire \sw_163_module_data_in[7] ;
 wire \sw_163_module_data_out[0] ;
 wire \sw_163_module_data_out[1] ;
 wire \sw_163_module_data_out[2] ;
 wire \sw_163_module_data_out[3] ;
 wire \sw_163_module_data_out[4] ;
 wire \sw_163_module_data_out[5] ;
 wire \sw_163_module_data_out[6] ;
 wire \sw_163_module_data_out[7] ;
 wire sw_163_scan_out;
 wire sw_164_clk_out;
 wire sw_164_data_out;
 wire sw_164_latch_out;
 wire \sw_164_module_data_in[0] ;
 wire \sw_164_module_data_in[1] ;
 wire \sw_164_module_data_in[2] ;
 wire \sw_164_module_data_in[3] ;
 wire \sw_164_module_data_in[4] ;
 wire \sw_164_module_data_in[5] ;
 wire \sw_164_module_data_in[6] ;
 wire \sw_164_module_data_in[7] ;
 wire \sw_164_module_data_out[0] ;
 wire \sw_164_module_data_out[1] ;
 wire \sw_164_module_data_out[2] ;
 wire \sw_164_module_data_out[3] ;
 wire \sw_164_module_data_out[4] ;
 wire \sw_164_module_data_out[5] ;
 wire \sw_164_module_data_out[6] ;
 wire \sw_164_module_data_out[7] ;
 wire sw_164_scan_out;
 wire sw_165_clk_out;
 wire sw_165_data_out;
 wire sw_165_latch_out;
 wire \sw_165_module_data_in[0] ;
 wire \sw_165_module_data_in[1] ;
 wire \sw_165_module_data_in[2] ;
 wire \sw_165_module_data_in[3] ;
 wire \sw_165_module_data_in[4] ;
 wire \sw_165_module_data_in[5] ;
 wire \sw_165_module_data_in[6] ;
 wire \sw_165_module_data_in[7] ;
 wire \sw_165_module_data_out[0] ;
 wire \sw_165_module_data_out[1] ;
 wire \sw_165_module_data_out[2] ;
 wire \sw_165_module_data_out[3] ;
 wire \sw_165_module_data_out[4] ;
 wire \sw_165_module_data_out[5] ;
 wire \sw_165_module_data_out[6] ;
 wire \sw_165_module_data_out[7] ;
 wire sw_165_scan_out;
 wire sw_166_clk_out;
 wire sw_166_data_out;
 wire sw_166_latch_out;
 wire \sw_166_module_data_in[0] ;
 wire \sw_166_module_data_in[1] ;
 wire \sw_166_module_data_in[2] ;
 wire \sw_166_module_data_in[3] ;
 wire \sw_166_module_data_in[4] ;
 wire \sw_166_module_data_in[5] ;
 wire \sw_166_module_data_in[6] ;
 wire \sw_166_module_data_in[7] ;
 wire \sw_166_module_data_out[0] ;
 wire \sw_166_module_data_out[1] ;
 wire \sw_166_module_data_out[2] ;
 wire \sw_166_module_data_out[3] ;
 wire \sw_166_module_data_out[4] ;
 wire \sw_166_module_data_out[5] ;
 wire \sw_166_module_data_out[6] ;
 wire \sw_166_module_data_out[7] ;
 wire sw_166_scan_out;
 wire sw_167_clk_out;
 wire sw_167_data_out;
 wire sw_167_latch_out;
 wire \sw_167_module_data_in[0] ;
 wire \sw_167_module_data_in[1] ;
 wire \sw_167_module_data_in[2] ;
 wire \sw_167_module_data_in[3] ;
 wire \sw_167_module_data_in[4] ;
 wire \sw_167_module_data_in[5] ;
 wire \sw_167_module_data_in[6] ;
 wire \sw_167_module_data_in[7] ;
 wire \sw_167_module_data_out[0] ;
 wire \sw_167_module_data_out[1] ;
 wire \sw_167_module_data_out[2] ;
 wire \sw_167_module_data_out[3] ;
 wire \sw_167_module_data_out[4] ;
 wire \sw_167_module_data_out[5] ;
 wire \sw_167_module_data_out[6] ;
 wire \sw_167_module_data_out[7] ;
 wire sw_167_scan_out;
 wire sw_168_clk_out;
 wire sw_168_data_out;
 wire sw_168_latch_out;
 wire \sw_168_module_data_in[0] ;
 wire \sw_168_module_data_in[1] ;
 wire \sw_168_module_data_in[2] ;
 wire \sw_168_module_data_in[3] ;
 wire \sw_168_module_data_in[4] ;
 wire \sw_168_module_data_in[5] ;
 wire \sw_168_module_data_in[6] ;
 wire \sw_168_module_data_in[7] ;
 wire \sw_168_module_data_out[0] ;
 wire \sw_168_module_data_out[1] ;
 wire \sw_168_module_data_out[2] ;
 wire \sw_168_module_data_out[3] ;
 wire \sw_168_module_data_out[4] ;
 wire \sw_168_module_data_out[5] ;
 wire \sw_168_module_data_out[6] ;
 wire \sw_168_module_data_out[7] ;
 wire sw_168_scan_out;
 wire sw_169_clk_out;
 wire sw_169_data_out;
 wire sw_169_latch_out;
 wire \sw_169_module_data_in[0] ;
 wire \sw_169_module_data_in[1] ;
 wire \sw_169_module_data_in[2] ;
 wire \sw_169_module_data_in[3] ;
 wire \sw_169_module_data_in[4] ;
 wire \sw_169_module_data_in[5] ;
 wire \sw_169_module_data_in[6] ;
 wire \sw_169_module_data_in[7] ;
 wire \sw_169_module_data_out[0] ;
 wire \sw_169_module_data_out[1] ;
 wire \sw_169_module_data_out[2] ;
 wire \sw_169_module_data_out[3] ;
 wire \sw_169_module_data_out[4] ;
 wire \sw_169_module_data_out[5] ;
 wire \sw_169_module_data_out[6] ;
 wire \sw_169_module_data_out[7] ;
 wire sw_169_scan_out;
 wire sw_170_clk_out;
 wire sw_170_data_out;
 wire sw_170_latch_out;
 wire \sw_170_module_data_in[0] ;
 wire \sw_170_module_data_in[1] ;
 wire \sw_170_module_data_in[2] ;
 wire \sw_170_module_data_in[3] ;
 wire \sw_170_module_data_in[4] ;
 wire \sw_170_module_data_in[5] ;
 wire \sw_170_module_data_in[6] ;
 wire \sw_170_module_data_in[7] ;
 wire \sw_170_module_data_out[0] ;
 wire \sw_170_module_data_out[1] ;
 wire \sw_170_module_data_out[2] ;
 wire \sw_170_module_data_out[3] ;
 wire \sw_170_module_data_out[4] ;
 wire \sw_170_module_data_out[5] ;
 wire \sw_170_module_data_out[6] ;
 wire \sw_170_module_data_out[7] ;
 wire sw_170_scan_out;
 wire sw_171_clk_out;
 wire sw_171_data_out;
 wire sw_171_latch_out;
 wire \sw_171_module_data_in[0] ;
 wire \sw_171_module_data_in[1] ;
 wire \sw_171_module_data_in[2] ;
 wire \sw_171_module_data_in[3] ;
 wire \sw_171_module_data_in[4] ;
 wire \sw_171_module_data_in[5] ;
 wire \sw_171_module_data_in[6] ;
 wire \sw_171_module_data_in[7] ;
 wire \sw_171_module_data_out[0] ;
 wire \sw_171_module_data_out[1] ;
 wire \sw_171_module_data_out[2] ;
 wire \sw_171_module_data_out[3] ;
 wire \sw_171_module_data_out[4] ;
 wire \sw_171_module_data_out[5] ;
 wire \sw_171_module_data_out[6] ;
 wire \sw_171_module_data_out[7] ;
 wire sw_171_scan_out;
 wire sw_172_clk_out;
 wire sw_172_data_out;
 wire sw_172_latch_out;
 wire \sw_172_module_data_in[0] ;
 wire \sw_172_module_data_in[1] ;
 wire \sw_172_module_data_in[2] ;
 wire \sw_172_module_data_in[3] ;
 wire \sw_172_module_data_in[4] ;
 wire \sw_172_module_data_in[5] ;
 wire \sw_172_module_data_in[6] ;
 wire \sw_172_module_data_in[7] ;
 wire \sw_172_module_data_out[0] ;
 wire \sw_172_module_data_out[1] ;
 wire \sw_172_module_data_out[2] ;
 wire \sw_172_module_data_out[3] ;
 wire \sw_172_module_data_out[4] ;
 wire \sw_172_module_data_out[5] ;
 wire \sw_172_module_data_out[6] ;
 wire \sw_172_module_data_out[7] ;
 wire sw_172_scan_out;
 wire sw_173_clk_out;
 wire sw_173_data_out;
 wire sw_173_latch_out;
 wire \sw_173_module_data_in[0] ;
 wire \sw_173_module_data_in[1] ;
 wire \sw_173_module_data_in[2] ;
 wire \sw_173_module_data_in[3] ;
 wire \sw_173_module_data_in[4] ;
 wire \sw_173_module_data_in[5] ;
 wire \sw_173_module_data_in[6] ;
 wire \sw_173_module_data_in[7] ;
 wire \sw_173_module_data_out[0] ;
 wire \sw_173_module_data_out[1] ;
 wire \sw_173_module_data_out[2] ;
 wire \sw_173_module_data_out[3] ;
 wire \sw_173_module_data_out[4] ;
 wire \sw_173_module_data_out[5] ;
 wire \sw_173_module_data_out[6] ;
 wire \sw_173_module_data_out[7] ;
 wire sw_173_scan_out;
 wire sw_174_clk_out;
 wire sw_174_data_out;
 wire sw_174_latch_out;
 wire \sw_174_module_data_in[0] ;
 wire \sw_174_module_data_in[1] ;
 wire \sw_174_module_data_in[2] ;
 wire \sw_174_module_data_in[3] ;
 wire \sw_174_module_data_in[4] ;
 wire \sw_174_module_data_in[5] ;
 wire \sw_174_module_data_in[6] ;
 wire \sw_174_module_data_in[7] ;
 wire \sw_174_module_data_out[0] ;
 wire \sw_174_module_data_out[1] ;
 wire \sw_174_module_data_out[2] ;
 wire \sw_174_module_data_out[3] ;
 wire \sw_174_module_data_out[4] ;
 wire \sw_174_module_data_out[5] ;
 wire \sw_174_module_data_out[6] ;
 wire \sw_174_module_data_out[7] ;
 wire sw_174_scan_out;
 wire sw_175_clk_out;
 wire sw_175_data_out;
 wire sw_175_latch_out;
 wire \sw_175_module_data_in[0] ;
 wire \sw_175_module_data_in[1] ;
 wire \sw_175_module_data_in[2] ;
 wire \sw_175_module_data_in[3] ;
 wire \sw_175_module_data_in[4] ;
 wire \sw_175_module_data_in[5] ;
 wire \sw_175_module_data_in[6] ;
 wire \sw_175_module_data_in[7] ;
 wire \sw_175_module_data_out[0] ;
 wire \sw_175_module_data_out[1] ;
 wire \sw_175_module_data_out[2] ;
 wire \sw_175_module_data_out[3] ;
 wire \sw_175_module_data_out[4] ;
 wire \sw_175_module_data_out[5] ;
 wire \sw_175_module_data_out[6] ;
 wire \sw_175_module_data_out[7] ;
 wire sw_175_scan_out;
 wire sw_176_clk_out;
 wire sw_176_data_out;
 wire sw_176_latch_out;
 wire \sw_176_module_data_in[0] ;
 wire \sw_176_module_data_in[1] ;
 wire \sw_176_module_data_in[2] ;
 wire \sw_176_module_data_in[3] ;
 wire \sw_176_module_data_in[4] ;
 wire \sw_176_module_data_in[5] ;
 wire \sw_176_module_data_in[6] ;
 wire \sw_176_module_data_in[7] ;
 wire \sw_176_module_data_out[0] ;
 wire \sw_176_module_data_out[1] ;
 wire \sw_176_module_data_out[2] ;
 wire \sw_176_module_data_out[3] ;
 wire \sw_176_module_data_out[4] ;
 wire \sw_176_module_data_out[5] ;
 wire \sw_176_module_data_out[6] ;
 wire \sw_176_module_data_out[7] ;
 wire sw_176_scan_out;
 wire sw_177_clk_out;
 wire sw_177_data_out;
 wire sw_177_latch_out;
 wire \sw_177_module_data_in[0] ;
 wire \sw_177_module_data_in[1] ;
 wire \sw_177_module_data_in[2] ;
 wire \sw_177_module_data_in[3] ;
 wire \sw_177_module_data_in[4] ;
 wire \sw_177_module_data_in[5] ;
 wire \sw_177_module_data_in[6] ;
 wire \sw_177_module_data_in[7] ;
 wire \sw_177_module_data_out[0] ;
 wire \sw_177_module_data_out[1] ;
 wire \sw_177_module_data_out[2] ;
 wire \sw_177_module_data_out[3] ;
 wire \sw_177_module_data_out[4] ;
 wire \sw_177_module_data_out[5] ;
 wire \sw_177_module_data_out[6] ;
 wire \sw_177_module_data_out[7] ;
 wire sw_177_scan_out;
 wire sw_178_clk_out;
 wire sw_178_data_out;
 wire sw_178_latch_out;
 wire \sw_178_module_data_in[0] ;
 wire \sw_178_module_data_in[1] ;
 wire \sw_178_module_data_in[2] ;
 wire \sw_178_module_data_in[3] ;
 wire \sw_178_module_data_in[4] ;
 wire \sw_178_module_data_in[5] ;
 wire \sw_178_module_data_in[6] ;
 wire \sw_178_module_data_in[7] ;
 wire \sw_178_module_data_out[0] ;
 wire \sw_178_module_data_out[1] ;
 wire \sw_178_module_data_out[2] ;
 wire \sw_178_module_data_out[3] ;
 wire \sw_178_module_data_out[4] ;
 wire \sw_178_module_data_out[5] ;
 wire \sw_178_module_data_out[6] ;
 wire \sw_178_module_data_out[7] ;
 wire sw_178_scan_out;
 wire sw_179_clk_out;
 wire sw_179_data_out;
 wire sw_179_latch_out;
 wire \sw_179_module_data_in[0] ;
 wire \sw_179_module_data_in[1] ;
 wire \sw_179_module_data_in[2] ;
 wire \sw_179_module_data_in[3] ;
 wire \sw_179_module_data_in[4] ;
 wire \sw_179_module_data_in[5] ;
 wire \sw_179_module_data_in[6] ;
 wire \sw_179_module_data_in[7] ;
 wire \sw_179_module_data_out[0] ;
 wire \sw_179_module_data_out[1] ;
 wire \sw_179_module_data_out[2] ;
 wire \sw_179_module_data_out[3] ;
 wire \sw_179_module_data_out[4] ;
 wire \sw_179_module_data_out[5] ;
 wire \sw_179_module_data_out[6] ;
 wire \sw_179_module_data_out[7] ;
 wire sw_179_scan_out;
 wire sw_180_clk_out;
 wire sw_180_data_out;
 wire sw_180_latch_out;
 wire \sw_180_module_data_in[0] ;
 wire \sw_180_module_data_in[1] ;
 wire \sw_180_module_data_in[2] ;
 wire \sw_180_module_data_in[3] ;
 wire \sw_180_module_data_in[4] ;
 wire \sw_180_module_data_in[5] ;
 wire \sw_180_module_data_in[6] ;
 wire \sw_180_module_data_in[7] ;
 wire \sw_180_module_data_out[0] ;
 wire \sw_180_module_data_out[1] ;
 wire \sw_180_module_data_out[2] ;
 wire \sw_180_module_data_out[3] ;
 wire \sw_180_module_data_out[4] ;
 wire \sw_180_module_data_out[5] ;
 wire \sw_180_module_data_out[6] ;
 wire \sw_180_module_data_out[7] ;
 wire sw_180_scan_out;
 wire sw_181_clk_out;
 wire sw_181_data_out;
 wire sw_181_latch_out;
 wire \sw_181_module_data_in[0] ;
 wire \sw_181_module_data_in[1] ;
 wire \sw_181_module_data_in[2] ;
 wire \sw_181_module_data_in[3] ;
 wire \sw_181_module_data_in[4] ;
 wire \sw_181_module_data_in[5] ;
 wire \sw_181_module_data_in[6] ;
 wire \sw_181_module_data_in[7] ;
 wire \sw_181_module_data_out[0] ;
 wire \sw_181_module_data_out[1] ;
 wire \sw_181_module_data_out[2] ;
 wire \sw_181_module_data_out[3] ;
 wire \sw_181_module_data_out[4] ;
 wire \sw_181_module_data_out[5] ;
 wire \sw_181_module_data_out[6] ;
 wire \sw_181_module_data_out[7] ;
 wire sw_181_scan_out;
 wire sw_182_clk_out;
 wire sw_182_data_out;
 wire sw_182_latch_out;
 wire \sw_182_module_data_in[0] ;
 wire \sw_182_module_data_in[1] ;
 wire \sw_182_module_data_in[2] ;
 wire \sw_182_module_data_in[3] ;
 wire \sw_182_module_data_in[4] ;
 wire \sw_182_module_data_in[5] ;
 wire \sw_182_module_data_in[6] ;
 wire \sw_182_module_data_in[7] ;
 wire \sw_182_module_data_out[0] ;
 wire \sw_182_module_data_out[1] ;
 wire \sw_182_module_data_out[2] ;
 wire \sw_182_module_data_out[3] ;
 wire \sw_182_module_data_out[4] ;
 wire \sw_182_module_data_out[5] ;
 wire \sw_182_module_data_out[6] ;
 wire \sw_182_module_data_out[7] ;
 wire sw_182_scan_out;
 wire sw_183_clk_out;
 wire sw_183_data_out;
 wire sw_183_latch_out;
 wire \sw_183_module_data_in[0] ;
 wire \sw_183_module_data_in[1] ;
 wire \sw_183_module_data_in[2] ;
 wire \sw_183_module_data_in[3] ;
 wire \sw_183_module_data_in[4] ;
 wire \sw_183_module_data_in[5] ;
 wire \sw_183_module_data_in[6] ;
 wire \sw_183_module_data_in[7] ;
 wire \sw_183_module_data_out[0] ;
 wire \sw_183_module_data_out[1] ;
 wire \sw_183_module_data_out[2] ;
 wire \sw_183_module_data_out[3] ;
 wire \sw_183_module_data_out[4] ;
 wire \sw_183_module_data_out[5] ;
 wire \sw_183_module_data_out[6] ;
 wire \sw_183_module_data_out[7] ;
 wire sw_183_scan_out;
 wire sw_184_clk_out;
 wire sw_184_data_out;
 wire sw_184_latch_out;
 wire \sw_184_module_data_in[0] ;
 wire \sw_184_module_data_in[1] ;
 wire \sw_184_module_data_in[2] ;
 wire \sw_184_module_data_in[3] ;
 wire \sw_184_module_data_in[4] ;
 wire \sw_184_module_data_in[5] ;
 wire \sw_184_module_data_in[6] ;
 wire \sw_184_module_data_in[7] ;
 wire \sw_184_module_data_out[0] ;
 wire \sw_184_module_data_out[1] ;
 wire \sw_184_module_data_out[2] ;
 wire \sw_184_module_data_out[3] ;
 wire \sw_184_module_data_out[4] ;
 wire \sw_184_module_data_out[5] ;
 wire \sw_184_module_data_out[6] ;
 wire \sw_184_module_data_out[7] ;
 wire sw_184_scan_out;
 wire sw_185_clk_out;
 wire sw_185_data_out;
 wire sw_185_latch_out;
 wire \sw_185_module_data_in[0] ;
 wire \sw_185_module_data_in[1] ;
 wire \sw_185_module_data_in[2] ;
 wire \sw_185_module_data_in[3] ;
 wire \sw_185_module_data_in[4] ;
 wire \sw_185_module_data_in[5] ;
 wire \sw_185_module_data_in[6] ;
 wire \sw_185_module_data_in[7] ;
 wire \sw_185_module_data_out[0] ;
 wire \sw_185_module_data_out[1] ;
 wire \sw_185_module_data_out[2] ;
 wire \sw_185_module_data_out[3] ;
 wire \sw_185_module_data_out[4] ;
 wire \sw_185_module_data_out[5] ;
 wire \sw_185_module_data_out[6] ;
 wire \sw_185_module_data_out[7] ;
 wire sw_185_scan_out;
 wire sw_186_clk_out;
 wire sw_186_data_out;
 wire sw_186_latch_out;
 wire \sw_186_module_data_in[0] ;
 wire \sw_186_module_data_in[1] ;
 wire \sw_186_module_data_in[2] ;
 wire \sw_186_module_data_in[3] ;
 wire \sw_186_module_data_in[4] ;
 wire \sw_186_module_data_in[5] ;
 wire \sw_186_module_data_in[6] ;
 wire \sw_186_module_data_in[7] ;
 wire \sw_186_module_data_out[0] ;
 wire \sw_186_module_data_out[1] ;
 wire \sw_186_module_data_out[2] ;
 wire \sw_186_module_data_out[3] ;
 wire \sw_186_module_data_out[4] ;
 wire \sw_186_module_data_out[5] ;
 wire \sw_186_module_data_out[6] ;
 wire \sw_186_module_data_out[7] ;
 wire sw_186_scan_out;
 wire sw_187_clk_out;
 wire sw_187_data_out;
 wire sw_187_latch_out;
 wire \sw_187_module_data_in[0] ;
 wire \sw_187_module_data_in[1] ;
 wire \sw_187_module_data_in[2] ;
 wire \sw_187_module_data_in[3] ;
 wire \sw_187_module_data_in[4] ;
 wire \sw_187_module_data_in[5] ;
 wire \sw_187_module_data_in[6] ;
 wire \sw_187_module_data_in[7] ;
 wire \sw_187_module_data_out[0] ;
 wire \sw_187_module_data_out[1] ;
 wire \sw_187_module_data_out[2] ;
 wire \sw_187_module_data_out[3] ;
 wire \sw_187_module_data_out[4] ;
 wire \sw_187_module_data_out[5] ;
 wire \sw_187_module_data_out[6] ;
 wire \sw_187_module_data_out[7] ;
 wire sw_187_scan_out;
 wire sw_188_clk_out;
 wire sw_188_data_out;
 wire sw_188_latch_out;
 wire \sw_188_module_data_in[0] ;
 wire \sw_188_module_data_in[1] ;
 wire \sw_188_module_data_in[2] ;
 wire \sw_188_module_data_in[3] ;
 wire \sw_188_module_data_in[4] ;
 wire \sw_188_module_data_in[5] ;
 wire \sw_188_module_data_in[6] ;
 wire \sw_188_module_data_in[7] ;
 wire \sw_188_module_data_out[0] ;
 wire \sw_188_module_data_out[1] ;
 wire \sw_188_module_data_out[2] ;
 wire \sw_188_module_data_out[3] ;
 wire \sw_188_module_data_out[4] ;
 wire \sw_188_module_data_out[5] ;
 wire \sw_188_module_data_out[6] ;
 wire \sw_188_module_data_out[7] ;
 wire sw_188_scan_out;
 wire sw_189_clk_out;
 wire sw_189_data_out;
 wire sw_189_latch_out;
 wire \sw_189_module_data_in[0] ;
 wire \sw_189_module_data_in[1] ;
 wire \sw_189_module_data_in[2] ;
 wire \sw_189_module_data_in[3] ;
 wire \sw_189_module_data_in[4] ;
 wire \sw_189_module_data_in[5] ;
 wire \sw_189_module_data_in[6] ;
 wire \sw_189_module_data_in[7] ;
 wire \sw_189_module_data_out[0] ;
 wire \sw_189_module_data_out[1] ;
 wire \sw_189_module_data_out[2] ;
 wire \sw_189_module_data_out[3] ;
 wire \sw_189_module_data_out[4] ;
 wire \sw_189_module_data_out[5] ;
 wire \sw_189_module_data_out[6] ;
 wire \sw_189_module_data_out[7] ;
 wire sw_189_scan_out;
 wire sw_190_clk_out;
 wire sw_190_data_out;
 wire sw_190_latch_out;
 wire \sw_190_module_data_in[0] ;
 wire \sw_190_module_data_in[1] ;
 wire \sw_190_module_data_in[2] ;
 wire \sw_190_module_data_in[3] ;
 wire \sw_190_module_data_in[4] ;
 wire \sw_190_module_data_in[5] ;
 wire \sw_190_module_data_in[6] ;
 wire \sw_190_module_data_in[7] ;
 wire \sw_190_module_data_out[0] ;
 wire \sw_190_module_data_out[1] ;
 wire \sw_190_module_data_out[2] ;
 wire \sw_190_module_data_out[3] ;
 wire \sw_190_module_data_out[4] ;
 wire \sw_190_module_data_out[5] ;
 wire \sw_190_module_data_out[6] ;
 wire \sw_190_module_data_out[7] ;
 wire sw_190_scan_out;
 wire sw_191_clk_out;
 wire sw_191_data_out;
 wire sw_191_latch_out;
 wire \sw_191_module_data_in[0] ;
 wire \sw_191_module_data_in[1] ;
 wire \sw_191_module_data_in[2] ;
 wire \sw_191_module_data_in[3] ;
 wire \sw_191_module_data_in[4] ;
 wire \sw_191_module_data_in[5] ;
 wire \sw_191_module_data_in[6] ;
 wire \sw_191_module_data_in[7] ;
 wire \sw_191_module_data_out[0] ;
 wire \sw_191_module_data_out[1] ;
 wire \sw_191_module_data_out[2] ;
 wire \sw_191_module_data_out[3] ;
 wire \sw_191_module_data_out[4] ;
 wire \sw_191_module_data_out[5] ;
 wire \sw_191_module_data_out[6] ;
 wire \sw_191_module_data_out[7] ;
 wire sw_191_scan_out;
 wire sw_192_clk_out;
 wire sw_192_data_out;
 wire sw_192_latch_out;
 wire \sw_192_module_data_in[0] ;
 wire \sw_192_module_data_in[1] ;
 wire \sw_192_module_data_in[2] ;
 wire \sw_192_module_data_in[3] ;
 wire \sw_192_module_data_in[4] ;
 wire \sw_192_module_data_in[5] ;
 wire \sw_192_module_data_in[6] ;
 wire \sw_192_module_data_in[7] ;
 wire \sw_192_module_data_out[0] ;
 wire \sw_192_module_data_out[1] ;
 wire \sw_192_module_data_out[2] ;
 wire \sw_192_module_data_out[3] ;
 wire \sw_192_module_data_out[4] ;
 wire \sw_192_module_data_out[5] ;
 wire \sw_192_module_data_out[6] ;
 wire \sw_192_module_data_out[7] ;
 wire sw_192_scan_out;
 wire sw_193_clk_out;
 wire sw_193_data_out;
 wire sw_193_latch_out;
 wire \sw_193_module_data_in[0] ;
 wire \sw_193_module_data_in[1] ;
 wire \sw_193_module_data_in[2] ;
 wire \sw_193_module_data_in[3] ;
 wire \sw_193_module_data_in[4] ;
 wire \sw_193_module_data_in[5] ;
 wire \sw_193_module_data_in[6] ;
 wire \sw_193_module_data_in[7] ;
 wire \sw_193_module_data_out[0] ;
 wire \sw_193_module_data_out[1] ;
 wire \sw_193_module_data_out[2] ;
 wire \sw_193_module_data_out[3] ;
 wire \sw_193_module_data_out[4] ;
 wire \sw_193_module_data_out[5] ;
 wire \sw_193_module_data_out[6] ;
 wire \sw_193_module_data_out[7] ;
 wire sw_193_scan_out;
 wire sw_194_clk_out;
 wire sw_194_data_out;
 wire sw_194_latch_out;
 wire \sw_194_module_data_in[0] ;
 wire \sw_194_module_data_in[1] ;
 wire \sw_194_module_data_in[2] ;
 wire \sw_194_module_data_in[3] ;
 wire \sw_194_module_data_in[4] ;
 wire \sw_194_module_data_in[5] ;
 wire \sw_194_module_data_in[6] ;
 wire \sw_194_module_data_in[7] ;
 wire \sw_194_module_data_out[0] ;
 wire \sw_194_module_data_out[1] ;
 wire \sw_194_module_data_out[2] ;
 wire \sw_194_module_data_out[3] ;
 wire \sw_194_module_data_out[4] ;
 wire \sw_194_module_data_out[5] ;
 wire \sw_194_module_data_out[6] ;
 wire \sw_194_module_data_out[7] ;
 wire sw_194_scan_out;
 wire sw_195_clk_out;
 wire sw_195_data_out;
 wire sw_195_latch_out;
 wire \sw_195_module_data_in[0] ;
 wire \sw_195_module_data_in[1] ;
 wire \sw_195_module_data_in[2] ;
 wire \sw_195_module_data_in[3] ;
 wire \sw_195_module_data_in[4] ;
 wire \sw_195_module_data_in[5] ;
 wire \sw_195_module_data_in[6] ;
 wire \sw_195_module_data_in[7] ;
 wire \sw_195_module_data_out[0] ;
 wire \sw_195_module_data_out[1] ;
 wire \sw_195_module_data_out[2] ;
 wire \sw_195_module_data_out[3] ;
 wire \sw_195_module_data_out[4] ;
 wire \sw_195_module_data_out[5] ;
 wire \sw_195_module_data_out[6] ;
 wire \sw_195_module_data_out[7] ;
 wire sw_195_scan_out;
 wire sw_196_clk_out;
 wire sw_196_data_out;
 wire sw_196_latch_out;
 wire \sw_196_module_data_in[0] ;
 wire \sw_196_module_data_in[1] ;
 wire \sw_196_module_data_in[2] ;
 wire \sw_196_module_data_in[3] ;
 wire \sw_196_module_data_in[4] ;
 wire \sw_196_module_data_in[5] ;
 wire \sw_196_module_data_in[6] ;
 wire \sw_196_module_data_in[7] ;
 wire \sw_196_module_data_out[0] ;
 wire \sw_196_module_data_out[1] ;
 wire \sw_196_module_data_out[2] ;
 wire \sw_196_module_data_out[3] ;
 wire \sw_196_module_data_out[4] ;
 wire \sw_196_module_data_out[5] ;
 wire \sw_196_module_data_out[6] ;
 wire \sw_196_module_data_out[7] ;
 wire sw_196_scan_out;
 wire sw_197_clk_out;
 wire sw_197_data_out;
 wire sw_197_latch_out;
 wire \sw_197_module_data_in[0] ;
 wire \sw_197_module_data_in[1] ;
 wire \sw_197_module_data_in[2] ;
 wire \sw_197_module_data_in[3] ;
 wire \sw_197_module_data_in[4] ;
 wire \sw_197_module_data_in[5] ;
 wire \sw_197_module_data_in[6] ;
 wire \sw_197_module_data_in[7] ;
 wire \sw_197_module_data_out[0] ;
 wire \sw_197_module_data_out[1] ;
 wire \sw_197_module_data_out[2] ;
 wire \sw_197_module_data_out[3] ;
 wire \sw_197_module_data_out[4] ;
 wire \sw_197_module_data_out[5] ;
 wire \sw_197_module_data_out[6] ;
 wire \sw_197_module_data_out[7] ;
 wire sw_197_scan_out;
 wire sw_198_clk_out;
 wire sw_198_data_out;
 wire sw_198_latch_out;
 wire \sw_198_module_data_in[0] ;
 wire \sw_198_module_data_in[1] ;
 wire \sw_198_module_data_in[2] ;
 wire \sw_198_module_data_in[3] ;
 wire \sw_198_module_data_in[4] ;
 wire \sw_198_module_data_in[5] ;
 wire \sw_198_module_data_in[6] ;
 wire \sw_198_module_data_in[7] ;
 wire \sw_198_module_data_out[0] ;
 wire \sw_198_module_data_out[1] ;
 wire \sw_198_module_data_out[2] ;
 wire \sw_198_module_data_out[3] ;
 wire \sw_198_module_data_out[4] ;
 wire \sw_198_module_data_out[5] ;
 wire \sw_198_module_data_out[6] ;
 wire \sw_198_module_data_out[7] ;
 wire sw_198_scan_out;
 wire sw_199_clk_out;
 wire sw_199_data_out;
 wire sw_199_latch_out;
 wire \sw_199_module_data_in[0] ;
 wire \sw_199_module_data_in[1] ;
 wire \sw_199_module_data_in[2] ;
 wire \sw_199_module_data_in[3] ;
 wire \sw_199_module_data_in[4] ;
 wire \sw_199_module_data_in[5] ;
 wire \sw_199_module_data_in[6] ;
 wire \sw_199_module_data_in[7] ;
 wire \sw_199_module_data_out[0] ;
 wire \sw_199_module_data_out[1] ;
 wire \sw_199_module_data_out[2] ;
 wire \sw_199_module_data_out[3] ;
 wire \sw_199_module_data_out[4] ;
 wire \sw_199_module_data_out[5] ;
 wire \sw_199_module_data_out[6] ;
 wire \sw_199_module_data_out[7] ;
 wire sw_199_scan_out;
 wire sw_200_clk_out;
 wire sw_200_data_out;
 wire sw_200_latch_out;
 wire \sw_200_module_data_in[0] ;
 wire \sw_200_module_data_in[1] ;
 wire \sw_200_module_data_in[2] ;
 wire \sw_200_module_data_in[3] ;
 wire \sw_200_module_data_in[4] ;
 wire \sw_200_module_data_in[5] ;
 wire \sw_200_module_data_in[6] ;
 wire \sw_200_module_data_in[7] ;
 wire \sw_200_module_data_out[0] ;
 wire \sw_200_module_data_out[1] ;
 wire \sw_200_module_data_out[2] ;
 wire \sw_200_module_data_out[3] ;
 wire \sw_200_module_data_out[4] ;
 wire \sw_200_module_data_out[5] ;
 wire \sw_200_module_data_out[6] ;
 wire \sw_200_module_data_out[7] ;
 wire sw_200_scan_out;
 wire sw_201_clk_out;
 wire sw_201_data_out;
 wire sw_201_latch_out;
 wire \sw_201_module_data_in[0] ;
 wire \sw_201_module_data_in[1] ;
 wire \sw_201_module_data_in[2] ;
 wire \sw_201_module_data_in[3] ;
 wire \sw_201_module_data_in[4] ;
 wire \sw_201_module_data_in[5] ;
 wire \sw_201_module_data_in[6] ;
 wire \sw_201_module_data_in[7] ;
 wire \sw_201_module_data_out[0] ;
 wire \sw_201_module_data_out[1] ;
 wire \sw_201_module_data_out[2] ;
 wire \sw_201_module_data_out[3] ;
 wire \sw_201_module_data_out[4] ;
 wire \sw_201_module_data_out[5] ;
 wire \sw_201_module_data_out[6] ;
 wire \sw_201_module_data_out[7] ;
 wire sw_201_scan_out;
 wire sw_202_clk_out;
 wire sw_202_data_out;
 wire sw_202_latch_out;
 wire \sw_202_module_data_in[0] ;
 wire \sw_202_module_data_in[1] ;
 wire \sw_202_module_data_in[2] ;
 wire \sw_202_module_data_in[3] ;
 wire \sw_202_module_data_in[4] ;
 wire \sw_202_module_data_in[5] ;
 wire \sw_202_module_data_in[6] ;
 wire \sw_202_module_data_in[7] ;
 wire \sw_202_module_data_out[0] ;
 wire \sw_202_module_data_out[1] ;
 wire \sw_202_module_data_out[2] ;
 wire \sw_202_module_data_out[3] ;
 wire \sw_202_module_data_out[4] ;
 wire \sw_202_module_data_out[5] ;
 wire \sw_202_module_data_out[6] ;
 wire \sw_202_module_data_out[7] ;
 wire sw_202_scan_out;
 wire sw_203_clk_out;
 wire sw_203_data_out;
 wire sw_203_latch_out;
 wire \sw_203_module_data_in[0] ;
 wire \sw_203_module_data_in[1] ;
 wire \sw_203_module_data_in[2] ;
 wire \sw_203_module_data_in[3] ;
 wire \sw_203_module_data_in[4] ;
 wire \sw_203_module_data_in[5] ;
 wire \sw_203_module_data_in[6] ;
 wire \sw_203_module_data_in[7] ;
 wire \sw_203_module_data_out[0] ;
 wire \sw_203_module_data_out[1] ;
 wire \sw_203_module_data_out[2] ;
 wire \sw_203_module_data_out[3] ;
 wire \sw_203_module_data_out[4] ;
 wire \sw_203_module_data_out[5] ;
 wire \sw_203_module_data_out[6] ;
 wire \sw_203_module_data_out[7] ;
 wire sw_203_scan_out;
 wire sw_204_clk_out;
 wire sw_204_data_out;
 wire sw_204_latch_out;
 wire \sw_204_module_data_in[0] ;
 wire \sw_204_module_data_in[1] ;
 wire \sw_204_module_data_in[2] ;
 wire \sw_204_module_data_in[3] ;
 wire \sw_204_module_data_in[4] ;
 wire \sw_204_module_data_in[5] ;
 wire \sw_204_module_data_in[6] ;
 wire \sw_204_module_data_in[7] ;
 wire \sw_204_module_data_out[0] ;
 wire \sw_204_module_data_out[1] ;
 wire \sw_204_module_data_out[2] ;
 wire \sw_204_module_data_out[3] ;
 wire \sw_204_module_data_out[4] ;
 wire \sw_204_module_data_out[5] ;
 wire \sw_204_module_data_out[6] ;
 wire \sw_204_module_data_out[7] ;
 wire sw_204_scan_out;
 wire sw_205_clk_out;
 wire sw_205_data_out;
 wire sw_205_latch_out;
 wire \sw_205_module_data_in[0] ;
 wire \sw_205_module_data_in[1] ;
 wire \sw_205_module_data_in[2] ;
 wire \sw_205_module_data_in[3] ;
 wire \sw_205_module_data_in[4] ;
 wire \sw_205_module_data_in[5] ;
 wire \sw_205_module_data_in[6] ;
 wire \sw_205_module_data_in[7] ;
 wire \sw_205_module_data_out[0] ;
 wire \sw_205_module_data_out[1] ;
 wire \sw_205_module_data_out[2] ;
 wire \sw_205_module_data_out[3] ;
 wire \sw_205_module_data_out[4] ;
 wire \sw_205_module_data_out[5] ;
 wire \sw_205_module_data_out[6] ;
 wire \sw_205_module_data_out[7] ;
 wire sw_205_scan_out;
 wire sw_206_clk_out;
 wire sw_206_data_out;
 wire sw_206_latch_out;
 wire \sw_206_module_data_in[0] ;
 wire \sw_206_module_data_in[1] ;
 wire \sw_206_module_data_in[2] ;
 wire \sw_206_module_data_in[3] ;
 wire \sw_206_module_data_in[4] ;
 wire \sw_206_module_data_in[5] ;
 wire \sw_206_module_data_in[6] ;
 wire \sw_206_module_data_in[7] ;
 wire \sw_206_module_data_out[0] ;
 wire \sw_206_module_data_out[1] ;
 wire \sw_206_module_data_out[2] ;
 wire \sw_206_module_data_out[3] ;
 wire \sw_206_module_data_out[4] ;
 wire \sw_206_module_data_out[5] ;
 wire \sw_206_module_data_out[6] ;
 wire \sw_206_module_data_out[7] ;
 wire sw_206_scan_out;
 wire sw_207_clk_out;
 wire sw_207_data_out;
 wire sw_207_latch_out;
 wire \sw_207_module_data_in[0] ;
 wire \sw_207_module_data_in[1] ;
 wire \sw_207_module_data_in[2] ;
 wire \sw_207_module_data_in[3] ;
 wire \sw_207_module_data_in[4] ;
 wire \sw_207_module_data_in[5] ;
 wire \sw_207_module_data_in[6] ;
 wire \sw_207_module_data_in[7] ;
 wire \sw_207_module_data_out[0] ;
 wire \sw_207_module_data_out[1] ;
 wire \sw_207_module_data_out[2] ;
 wire \sw_207_module_data_out[3] ;
 wire \sw_207_module_data_out[4] ;
 wire \sw_207_module_data_out[5] ;
 wire \sw_207_module_data_out[6] ;
 wire \sw_207_module_data_out[7] ;
 wire sw_207_scan_out;
 wire sw_208_clk_out;
 wire sw_208_data_out;
 wire sw_208_latch_out;
 wire \sw_208_module_data_in[0] ;
 wire \sw_208_module_data_in[1] ;
 wire \sw_208_module_data_in[2] ;
 wire \sw_208_module_data_in[3] ;
 wire \sw_208_module_data_in[4] ;
 wire \sw_208_module_data_in[5] ;
 wire \sw_208_module_data_in[6] ;
 wire \sw_208_module_data_in[7] ;
 wire \sw_208_module_data_out[0] ;
 wire \sw_208_module_data_out[1] ;
 wire \sw_208_module_data_out[2] ;
 wire \sw_208_module_data_out[3] ;
 wire \sw_208_module_data_out[4] ;
 wire \sw_208_module_data_out[5] ;
 wire \sw_208_module_data_out[6] ;
 wire \sw_208_module_data_out[7] ;
 wire sw_208_scan_out;
 wire sw_209_clk_out;
 wire sw_209_data_out;
 wire sw_209_latch_out;
 wire \sw_209_module_data_in[0] ;
 wire \sw_209_module_data_in[1] ;
 wire \sw_209_module_data_in[2] ;
 wire \sw_209_module_data_in[3] ;
 wire \sw_209_module_data_in[4] ;
 wire \sw_209_module_data_in[5] ;
 wire \sw_209_module_data_in[6] ;
 wire \sw_209_module_data_in[7] ;
 wire \sw_209_module_data_out[0] ;
 wire \sw_209_module_data_out[1] ;
 wire \sw_209_module_data_out[2] ;
 wire \sw_209_module_data_out[3] ;
 wire \sw_209_module_data_out[4] ;
 wire \sw_209_module_data_out[5] ;
 wire \sw_209_module_data_out[6] ;
 wire \sw_209_module_data_out[7] ;
 wire sw_209_scan_out;
 wire sw_210_clk_out;
 wire sw_210_data_out;
 wire sw_210_latch_out;
 wire \sw_210_module_data_in[0] ;
 wire \sw_210_module_data_in[1] ;
 wire \sw_210_module_data_in[2] ;
 wire \sw_210_module_data_in[3] ;
 wire \sw_210_module_data_in[4] ;
 wire \sw_210_module_data_in[5] ;
 wire \sw_210_module_data_in[6] ;
 wire \sw_210_module_data_in[7] ;
 wire \sw_210_module_data_out[0] ;
 wire \sw_210_module_data_out[1] ;
 wire \sw_210_module_data_out[2] ;
 wire \sw_210_module_data_out[3] ;
 wire \sw_210_module_data_out[4] ;
 wire \sw_210_module_data_out[5] ;
 wire \sw_210_module_data_out[6] ;
 wire \sw_210_module_data_out[7] ;
 wire sw_210_scan_out;
 wire sw_211_clk_out;
 wire sw_211_data_out;
 wire sw_211_latch_out;
 wire \sw_211_module_data_in[0] ;
 wire \sw_211_module_data_in[1] ;
 wire \sw_211_module_data_in[2] ;
 wire \sw_211_module_data_in[3] ;
 wire \sw_211_module_data_in[4] ;
 wire \sw_211_module_data_in[5] ;
 wire \sw_211_module_data_in[6] ;
 wire \sw_211_module_data_in[7] ;
 wire \sw_211_module_data_out[0] ;
 wire \sw_211_module_data_out[1] ;
 wire \sw_211_module_data_out[2] ;
 wire \sw_211_module_data_out[3] ;
 wire \sw_211_module_data_out[4] ;
 wire \sw_211_module_data_out[5] ;
 wire \sw_211_module_data_out[6] ;
 wire \sw_211_module_data_out[7] ;
 wire sw_211_scan_out;
 wire sw_212_clk_out;
 wire sw_212_data_out;
 wire sw_212_latch_out;
 wire \sw_212_module_data_in[0] ;
 wire \sw_212_module_data_in[1] ;
 wire \sw_212_module_data_in[2] ;
 wire \sw_212_module_data_in[3] ;
 wire \sw_212_module_data_in[4] ;
 wire \sw_212_module_data_in[5] ;
 wire \sw_212_module_data_in[6] ;
 wire \sw_212_module_data_in[7] ;
 wire \sw_212_module_data_out[0] ;
 wire \sw_212_module_data_out[1] ;
 wire \sw_212_module_data_out[2] ;
 wire \sw_212_module_data_out[3] ;
 wire \sw_212_module_data_out[4] ;
 wire \sw_212_module_data_out[5] ;
 wire \sw_212_module_data_out[6] ;
 wire \sw_212_module_data_out[7] ;
 wire sw_212_scan_out;
 wire sw_213_clk_out;
 wire sw_213_data_out;
 wire sw_213_latch_out;
 wire \sw_213_module_data_in[0] ;
 wire \sw_213_module_data_in[1] ;
 wire \sw_213_module_data_in[2] ;
 wire \sw_213_module_data_in[3] ;
 wire \sw_213_module_data_in[4] ;
 wire \sw_213_module_data_in[5] ;
 wire \sw_213_module_data_in[6] ;
 wire \sw_213_module_data_in[7] ;
 wire \sw_213_module_data_out[0] ;
 wire \sw_213_module_data_out[1] ;
 wire \sw_213_module_data_out[2] ;
 wire \sw_213_module_data_out[3] ;
 wire \sw_213_module_data_out[4] ;
 wire \sw_213_module_data_out[5] ;
 wire \sw_213_module_data_out[6] ;
 wire \sw_213_module_data_out[7] ;
 wire sw_213_scan_out;
 wire sw_214_clk_out;
 wire sw_214_data_out;
 wire sw_214_latch_out;
 wire \sw_214_module_data_in[0] ;
 wire \sw_214_module_data_in[1] ;
 wire \sw_214_module_data_in[2] ;
 wire \sw_214_module_data_in[3] ;
 wire \sw_214_module_data_in[4] ;
 wire \sw_214_module_data_in[5] ;
 wire \sw_214_module_data_in[6] ;
 wire \sw_214_module_data_in[7] ;
 wire \sw_214_module_data_out[0] ;
 wire \sw_214_module_data_out[1] ;
 wire \sw_214_module_data_out[2] ;
 wire \sw_214_module_data_out[3] ;
 wire \sw_214_module_data_out[4] ;
 wire \sw_214_module_data_out[5] ;
 wire \sw_214_module_data_out[6] ;
 wire \sw_214_module_data_out[7] ;
 wire sw_214_scan_out;
 wire sw_215_clk_out;
 wire sw_215_data_out;
 wire sw_215_latch_out;
 wire \sw_215_module_data_in[0] ;
 wire \sw_215_module_data_in[1] ;
 wire \sw_215_module_data_in[2] ;
 wire \sw_215_module_data_in[3] ;
 wire \sw_215_module_data_in[4] ;
 wire \sw_215_module_data_in[5] ;
 wire \sw_215_module_data_in[6] ;
 wire \sw_215_module_data_in[7] ;
 wire \sw_215_module_data_out[0] ;
 wire \sw_215_module_data_out[1] ;
 wire \sw_215_module_data_out[2] ;
 wire \sw_215_module_data_out[3] ;
 wire \sw_215_module_data_out[4] ;
 wire \sw_215_module_data_out[5] ;
 wire \sw_215_module_data_out[6] ;
 wire \sw_215_module_data_out[7] ;
 wire sw_215_scan_out;
 wire sw_216_clk_out;
 wire sw_216_data_out;
 wire sw_216_latch_out;
 wire \sw_216_module_data_in[0] ;
 wire \sw_216_module_data_in[1] ;
 wire \sw_216_module_data_in[2] ;
 wire \sw_216_module_data_in[3] ;
 wire \sw_216_module_data_in[4] ;
 wire \sw_216_module_data_in[5] ;
 wire \sw_216_module_data_in[6] ;
 wire \sw_216_module_data_in[7] ;
 wire \sw_216_module_data_out[0] ;
 wire \sw_216_module_data_out[1] ;
 wire \sw_216_module_data_out[2] ;
 wire \sw_216_module_data_out[3] ;
 wire \sw_216_module_data_out[4] ;
 wire \sw_216_module_data_out[5] ;
 wire \sw_216_module_data_out[6] ;
 wire \sw_216_module_data_out[7] ;
 wire sw_216_scan_out;
 wire sw_217_clk_out;
 wire sw_217_data_out;
 wire sw_217_latch_out;
 wire \sw_217_module_data_in[0] ;
 wire \sw_217_module_data_in[1] ;
 wire \sw_217_module_data_in[2] ;
 wire \sw_217_module_data_in[3] ;
 wire \sw_217_module_data_in[4] ;
 wire \sw_217_module_data_in[5] ;
 wire \sw_217_module_data_in[6] ;
 wire \sw_217_module_data_in[7] ;
 wire \sw_217_module_data_out[0] ;
 wire \sw_217_module_data_out[1] ;
 wire \sw_217_module_data_out[2] ;
 wire \sw_217_module_data_out[3] ;
 wire \sw_217_module_data_out[4] ;
 wire \sw_217_module_data_out[5] ;
 wire \sw_217_module_data_out[6] ;
 wire \sw_217_module_data_out[7] ;
 wire sw_217_scan_out;
 wire sw_218_clk_out;
 wire sw_218_data_out;
 wire sw_218_latch_out;
 wire \sw_218_module_data_in[0] ;
 wire \sw_218_module_data_in[1] ;
 wire \sw_218_module_data_in[2] ;
 wire \sw_218_module_data_in[3] ;
 wire \sw_218_module_data_in[4] ;
 wire \sw_218_module_data_in[5] ;
 wire \sw_218_module_data_in[6] ;
 wire \sw_218_module_data_in[7] ;
 wire \sw_218_module_data_out[0] ;
 wire \sw_218_module_data_out[1] ;
 wire \sw_218_module_data_out[2] ;
 wire \sw_218_module_data_out[3] ;
 wire \sw_218_module_data_out[4] ;
 wire \sw_218_module_data_out[5] ;
 wire \sw_218_module_data_out[6] ;
 wire \sw_218_module_data_out[7] ;
 wire sw_218_scan_out;
 wire sw_219_clk_out;
 wire sw_219_data_out;
 wire sw_219_latch_out;
 wire \sw_219_module_data_in[0] ;
 wire \sw_219_module_data_in[1] ;
 wire \sw_219_module_data_in[2] ;
 wire \sw_219_module_data_in[3] ;
 wire \sw_219_module_data_in[4] ;
 wire \sw_219_module_data_in[5] ;
 wire \sw_219_module_data_in[6] ;
 wire \sw_219_module_data_in[7] ;
 wire \sw_219_module_data_out[0] ;
 wire \sw_219_module_data_out[1] ;
 wire \sw_219_module_data_out[2] ;
 wire \sw_219_module_data_out[3] ;
 wire \sw_219_module_data_out[4] ;
 wire \sw_219_module_data_out[5] ;
 wire \sw_219_module_data_out[6] ;
 wire \sw_219_module_data_out[7] ;
 wire sw_219_scan_out;
 wire sw_220_clk_out;
 wire sw_220_data_out;
 wire sw_220_latch_out;
 wire \sw_220_module_data_in[0] ;
 wire \sw_220_module_data_in[1] ;
 wire \sw_220_module_data_in[2] ;
 wire \sw_220_module_data_in[3] ;
 wire \sw_220_module_data_in[4] ;
 wire \sw_220_module_data_in[5] ;
 wire \sw_220_module_data_in[6] ;
 wire \sw_220_module_data_in[7] ;
 wire \sw_220_module_data_out[0] ;
 wire \sw_220_module_data_out[1] ;
 wire \sw_220_module_data_out[2] ;
 wire \sw_220_module_data_out[3] ;
 wire \sw_220_module_data_out[4] ;
 wire \sw_220_module_data_out[5] ;
 wire \sw_220_module_data_out[6] ;
 wire \sw_220_module_data_out[7] ;
 wire sw_220_scan_out;
 wire sw_221_clk_out;
 wire sw_221_data_out;
 wire sw_221_latch_out;
 wire \sw_221_module_data_in[0] ;
 wire \sw_221_module_data_in[1] ;
 wire \sw_221_module_data_in[2] ;
 wire \sw_221_module_data_in[3] ;
 wire \sw_221_module_data_in[4] ;
 wire \sw_221_module_data_in[5] ;
 wire \sw_221_module_data_in[6] ;
 wire \sw_221_module_data_in[7] ;
 wire \sw_221_module_data_out[0] ;
 wire \sw_221_module_data_out[1] ;
 wire \sw_221_module_data_out[2] ;
 wire \sw_221_module_data_out[3] ;
 wire \sw_221_module_data_out[4] ;
 wire \sw_221_module_data_out[5] ;
 wire \sw_221_module_data_out[6] ;
 wire \sw_221_module_data_out[7] ;
 wire sw_221_scan_out;
 wire sw_222_clk_out;
 wire sw_222_data_out;
 wire sw_222_latch_out;
 wire \sw_222_module_data_in[0] ;
 wire \sw_222_module_data_in[1] ;
 wire \sw_222_module_data_in[2] ;
 wire \sw_222_module_data_in[3] ;
 wire \sw_222_module_data_in[4] ;
 wire \sw_222_module_data_in[5] ;
 wire \sw_222_module_data_in[6] ;
 wire \sw_222_module_data_in[7] ;
 wire \sw_222_module_data_out[0] ;
 wire \sw_222_module_data_out[1] ;
 wire \sw_222_module_data_out[2] ;
 wire \sw_222_module_data_out[3] ;
 wire \sw_222_module_data_out[4] ;
 wire \sw_222_module_data_out[5] ;
 wire \sw_222_module_data_out[6] ;
 wire \sw_222_module_data_out[7] ;
 wire sw_222_scan_out;
 wire sw_223_clk_out;
 wire sw_223_data_out;
 wire sw_223_latch_out;
 wire \sw_223_module_data_in[0] ;
 wire \sw_223_module_data_in[1] ;
 wire \sw_223_module_data_in[2] ;
 wire \sw_223_module_data_in[3] ;
 wire \sw_223_module_data_in[4] ;
 wire \sw_223_module_data_in[5] ;
 wire \sw_223_module_data_in[6] ;
 wire \sw_223_module_data_in[7] ;
 wire \sw_223_module_data_out[0] ;
 wire \sw_223_module_data_out[1] ;
 wire \sw_223_module_data_out[2] ;
 wire \sw_223_module_data_out[3] ;
 wire \sw_223_module_data_out[4] ;
 wire \sw_223_module_data_out[5] ;
 wire \sw_223_module_data_out[6] ;
 wire \sw_223_module_data_out[7] ;
 wire sw_223_scan_out;
 wire sw_224_clk_out;
 wire sw_224_data_out;
 wire sw_224_latch_out;
 wire \sw_224_module_data_in[0] ;
 wire \sw_224_module_data_in[1] ;
 wire \sw_224_module_data_in[2] ;
 wire \sw_224_module_data_in[3] ;
 wire \sw_224_module_data_in[4] ;
 wire \sw_224_module_data_in[5] ;
 wire \sw_224_module_data_in[6] ;
 wire \sw_224_module_data_in[7] ;
 wire \sw_224_module_data_out[0] ;
 wire \sw_224_module_data_out[1] ;
 wire \sw_224_module_data_out[2] ;
 wire \sw_224_module_data_out[3] ;
 wire \sw_224_module_data_out[4] ;
 wire \sw_224_module_data_out[5] ;
 wire \sw_224_module_data_out[6] ;
 wire \sw_224_module_data_out[7] ;
 wire sw_224_scan_out;
 wire sw_225_clk_out;
 wire sw_225_data_out;
 wire sw_225_latch_out;
 wire \sw_225_module_data_in[0] ;
 wire \sw_225_module_data_in[1] ;
 wire \sw_225_module_data_in[2] ;
 wire \sw_225_module_data_in[3] ;
 wire \sw_225_module_data_in[4] ;
 wire \sw_225_module_data_in[5] ;
 wire \sw_225_module_data_in[6] ;
 wire \sw_225_module_data_in[7] ;
 wire \sw_225_module_data_out[0] ;
 wire \sw_225_module_data_out[1] ;
 wire \sw_225_module_data_out[2] ;
 wire \sw_225_module_data_out[3] ;
 wire \sw_225_module_data_out[4] ;
 wire \sw_225_module_data_out[5] ;
 wire \sw_225_module_data_out[6] ;
 wire \sw_225_module_data_out[7] ;
 wire sw_225_scan_out;
 wire sw_226_clk_out;
 wire sw_226_data_out;
 wire sw_226_latch_out;
 wire \sw_226_module_data_in[0] ;
 wire \sw_226_module_data_in[1] ;
 wire \sw_226_module_data_in[2] ;
 wire \sw_226_module_data_in[3] ;
 wire \sw_226_module_data_in[4] ;
 wire \sw_226_module_data_in[5] ;
 wire \sw_226_module_data_in[6] ;
 wire \sw_226_module_data_in[7] ;
 wire \sw_226_module_data_out[0] ;
 wire \sw_226_module_data_out[1] ;
 wire \sw_226_module_data_out[2] ;
 wire \sw_226_module_data_out[3] ;
 wire \sw_226_module_data_out[4] ;
 wire \sw_226_module_data_out[5] ;
 wire \sw_226_module_data_out[6] ;
 wire \sw_226_module_data_out[7] ;
 wire sw_226_scan_out;
 wire sw_227_clk_out;
 wire sw_227_data_out;
 wire sw_227_latch_out;
 wire \sw_227_module_data_in[0] ;
 wire \sw_227_module_data_in[1] ;
 wire \sw_227_module_data_in[2] ;
 wire \sw_227_module_data_in[3] ;
 wire \sw_227_module_data_in[4] ;
 wire \sw_227_module_data_in[5] ;
 wire \sw_227_module_data_in[6] ;
 wire \sw_227_module_data_in[7] ;
 wire \sw_227_module_data_out[0] ;
 wire \sw_227_module_data_out[1] ;
 wire \sw_227_module_data_out[2] ;
 wire \sw_227_module_data_out[3] ;
 wire \sw_227_module_data_out[4] ;
 wire \sw_227_module_data_out[5] ;
 wire \sw_227_module_data_out[6] ;
 wire \sw_227_module_data_out[7] ;
 wire sw_227_scan_out;
 wire sw_228_clk_out;
 wire sw_228_data_out;
 wire sw_228_latch_out;
 wire \sw_228_module_data_in[0] ;
 wire \sw_228_module_data_in[1] ;
 wire \sw_228_module_data_in[2] ;
 wire \sw_228_module_data_in[3] ;
 wire \sw_228_module_data_in[4] ;
 wire \sw_228_module_data_in[5] ;
 wire \sw_228_module_data_in[6] ;
 wire \sw_228_module_data_in[7] ;
 wire \sw_228_module_data_out[0] ;
 wire \sw_228_module_data_out[1] ;
 wire \sw_228_module_data_out[2] ;
 wire \sw_228_module_data_out[3] ;
 wire \sw_228_module_data_out[4] ;
 wire \sw_228_module_data_out[5] ;
 wire \sw_228_module_data_out[6] ;
 wire \sw_228_module_data_out[7] ;
 wire sw_228_scan_out;
 wire sw_229_clk_out;
 wire sw_229_data_out;
 wire sw_229_latch_out;
 wire \sw_229_module_data_in[0] ;
 wire \sw_229_module_data_in[1] ;
 wire \sw_229_module_data_in[2] ;
 wire \sw_229_module_data_in[3] ;
 wire \sw_229_module_data_in[4] ;
 wire \sw_229_module_data_in[5] ;
 wire \sw_229_module_data_in[6] ;
 wire \sw_229_module_data_in[7] ;
 wire \sw_229_module_data_out[0] ;
 wire \sw_229_module_data_out[1] ;
 wire \sw_229_module_data_out[2] ;
 wire \sw_229_module_data_out[3] ;
 wire \sw_229_module_data_out[4] ;
 wire \sw_229_module_data_out[5] ;
 wire \sw_229_module_data_out[6] ;
 wire \sw_229_module_data_out[7] ;
 wire sw_229_scan_out;
 wire sw_230_clk_out;
 wire sw_230_data_out;
 wire sw_230_latch_out;
 wire \sw_230_module_data_in[0] ;
 wire \sw_230_module_data_in[1] ;
 wire \sw_230_module_data_in[2] ;
 wire \sw_230_module_data_in[3] ;
 wire \sw_230_module_data_in[4] ;
 wire \sw_230_module_data_in[5] ;
 wire \sw_230_module_data_in[6] ;
 wire \sw_230_module_data_in[7] ;
 wire \sw_230_module_data_out[0] ;
 wire \sw_230_module_data_out[1] ;
 wire \sw_230_module_data_out[2] ;
 wire \sw_230_module_data_out[3] ;
 wire \sw_230_module_data_out[4] ;
 wire \sw_230_module_data_out[5] ;
 wire \sw_230_module_data_out[6] ;
 wire \sw_230_module_data_out[7] ;
 wire sw_230_scan_out;
 wire sw_231_clk_out;
 wire sw_231_data_out;
 wire sw_231_latch_out;
 wire \sw_231_module_data_in[0] ;
 wire \sw_231_module_data_in[1] ;
 wire \sw_231_module_data_in[2] ;
 wire \sw_231_module_data_in[3] ;
 wire \sw_231_module_data_in[4] ;
 wire \sw_231_module_data_in[5] ;
 wire \sw_231_module_data_in[6] ;
 wire \sw_231_module_data_in[7] ;
 wire \sw_231_module_data_out[0] ;
 wire \sw_231_module_data_out[1] ;
 wire \sw_231_module_data_out[2] ;
 wire \sw_231_module_data_out[3] ;
 wire \sw_231_module_data_out[4] ;
 wire \sw_231_module_data_out[5] ;
 wire \sw_231_module_data_out[6] ;
 wire \sw_231_module_data_out[7] ;
 wire sw_231_scan_out;
 wire sw_232_clk_out;
 wire sw_232_data_out;
 wire sw_232_latch_out;
 wire \sw_232_module_data_in[0] ;
 wire \sw_232_module_data_in[1] ;
 wire \sw_232_module_data_in[2] ;
 wire \sw_232_module_data_in[3] ;
 wire \sw_232_module_data_in[4] ;
 wire \sw_232_module_data_in[5] ;
 wire \sw_232_module_data_in[6] ;
 wire \sw_232_module_data_in[7] ;
 wire \sw_232_module_data_out[0] ;
 wire \sw_232_module_data_out[1] ;
 wire \sw_232_module_data_out[2] ;
 wire \sw_232_module_data_out[3] ;
 wire \sw_232_module_data_out[4] ;
 wire \sw_232_module_data_out[5] ;
 wire \sw_232_module_data_out[6] ;
 wire \sw_232_module_data_out[7] ;
 wire sw_232_scan_out;
 wire sw_233_clk_out;
 wire sw_233_data_out;
 wire sw_233_latch_out;
 wire \sw_233_module_data_in[0] ;
 wire \sw_233_module_data_in[1] ;
 wire \sw_233_module_data_in[2] ;
 wire \sw_233_module_data_in[3] ;
 wire \sw_233_module_data_in[4] ;
 wire \sw_233_module_data_in[5] ;
 wire \sw_233_module_data_in[6] ;
 wire \sw_233_module_data_in[7] ;
 wire \sw_233_module_data_out[0] ;
 wire \sw_233_module_data_out[1] ;
 wire \sw_233_module_data_out[2] ;
 wire \sw_233_module_data_out[3] ;
 wire \sw_233_module_data_out[4] ;
 wire \sw_233_module_data_out[5] ;
 wire \sw_233_module_data_out[6] ;
 wire \sw_233_module_data_out[7] ;
 wire sw_233_scan_out;
 wire sw_234_clk_out;
 wire sw_234_data_out;
 wire sw_234_latch_out;
 wire \sw_234_module_data_in[0] ;
 wire \sw_234_module_data_in[1] ;
 wire \sw_234_module_data_in[2] ;
 wire \sw_234_module_data_in[3] ;
 wire \sw_234_module_data_in[4] ;
 wire \sw_234_module_data_in[5] ;
 wire \sw_234_module_data_in[6] ;
 wire \sw_234_module_data_in[7] ;
 wire \sw_234_module_data_out[0] ;
 wire \sw_234_module_data_out[1] ;
 wire \sw_234_module_data_out[2] ;
 wire \sw_234_module_data_out[3] ;
 wire \sw_234_module_data_out[4] ;
 wire \sw_234_module_data_out[5] ;
 wire \sw_234_module_data_out[6] ;
 wire \sw_234_module_data_out[7] ;
 wire sw_234_scan_out;
 wire sw_235_clk_out;
 wire sw_235_data_out;
 wire sw_235_latch_out;
 wire \sw_235_module_data_in[0] ;
 wire \sw_235_module_data_in[1] ;
 wire \sw_235_module_data_in[2] ;
 wire \sw_235_module_data_in[3] ;
 wire \sw_235_module_data_in[4] ;
 wire \sw_235_module_data_in[5] ;
 wire \sw_235_module_data_in[6] ;
 wire \sw_235_module_data_in[7] ;
 wire \sw_235_module_data_out[0] ;
 wire \sw_235_module_data_out[1] ;
 wire \sw_235_module_data_out[2] ;
 wire \sw_235_module_data_out[3] ;
 wire \sw_235_module_data_out[4] ;
 wire \sw_235_module_data_out[5] ;
 wire \sw_235_module_data_out[6] ;
 wire \sw_235_module_data_out[7] ;
 wire sw_235_scan_out;
 wire sw_236_clk_out;
 wire sw_236_data_out;
 wire sw_236_latch_out;
 wire \sw_236_module_data_in[0] ;
 wire \sw_236_module_data_in[1] ;
 wire \sw_236_module_data_in[2] ;
 wire \sw_236_module_data_in[3] ;
 wire \sw_236_module_data_in[4] ;
 wire \sw_236_module_data_in[5] ;
 wire \sw_236_module_data_in[6] ;
 wire \sw_236_module_data_in[7] ;
 wire \sw_236_module_data_out[0] ;
 wire \sw_236_module_data_out[1] ;
 wire \sw_236_module_data_out[2] ;
 wire \sw_236_module_data_out[3] ;
 wire \sw_236_module_data_out[4] ;
 wire \sw_236_module_data_out[5] ;
 wire \sw_236_module_data_out[6] ;
 wire \sw_236_module_data_out[7] ;
 wire sw_236_scan_out;
 wire sw_237_clk_out;
 wire sw_237_data_out;
 wire sw_237_latch_out;
 wire \sw_237_module_data_in[0] ;
 wire \sw_237_module_data_in[1] ;
 wire \sw_237_module_data_in[2] ;
 wire \sw_237_module_data_in[3] ;
 wire \sw_237_module_data_in[4] ;
 wire \sw_237_module_data_in[5] ;
 wire \sw_237_module_data_in[6] ;
 wire \sw_237_module_data_in[7] ;
 wire \sw_237_module_data_out[0] ;
 wire \sw_237_module_data_out[1] ;
 wire \sw_237_module_data_out[2] ;
 wire \sw_237_module_data_out[3] ;
 wire \sw_237_module_data_out[4] ;
 wire \sw_237_module_data_out[5] ;
 wire \sw_237_module_data_out[6] ;
 wire \sw_237_module_data_out[7] ;
 wire sw_237_scan_out;
 wire sw_238_clk_out;
 wire sw_238_data_out;
 wire sw_238_latch_out;
 wire \sw_238_module_data_in[0] ;
 wire \sw_238_module_data_in[1] ;
 wire \sw_238_module_data_in[2] ;
 wire \sw_238_module_data_in[3] ;
 wire \sw_238_module_data_in[4] ;
 wire \sw_238_module_data_in[5] ;
 wire \sw_238_module_data_in[6] ;
 wire \sw_238_module_data_in[7] ;
 wire \sw_238_module_data_out[0] ;
 wire \sw_238_module_data_out[1] ;
 wire \sw_238_module_data_out[2] ;
 wire \sw_238_module_data_out[3] ;
 wire \sw_238_module_data_out[4] ;
 wire \sw_238_module_data_out[5] ;
 wire \sw_238_module_data_out[6] ;
 wire \sw_238_module_data_out[7] ;
 wire sw_238_scan_out;
 wire sw_239_clk_out;
 wire sw_239_data_out;
 wire sw_239_latch_out;
 wire \sw_239_module_data_in[0] ;
 wire \sw_239_module_data_in[1] ;
 wire \sw_239_module_data_in[2] ;
 wire \sw_239_module_data_in[3] ;
 wire \sw_239_module_data_in[4] ;
 wire \sw_239_module_data_in[5] ;
 wire \sw_239_module_data_in[6] ;
 wire \sw_239_module_data_in[7] ;
 wire \sw_239_module_data_out[0] ;
 wire \sw_239_module_data_out[1] ;
 wire \sw_239_module_data_out[2] ;
 wire \sw_239_module_data_out[3] ;
 wire \sw_239_module_data_out[4] ;
 wire \sw_239_module_data_out[5] ;
 wire \sw_239_module_data_out[6] ;
 wire \sw_239_module_data_out[7] ;
 wire sw_239_scan_out;
 wire sw_240_clk_out;
 wire sw_240_data_out;
 wire sw_240_latch_out;
 wire \sw_240_module_data_in[0] ;
 wire \sw_240_module_data_in[1] ;
 wire \sw_240_module_data_in[2] ;
 wire \sw_240_module_data_in[3] ;
 wire \sw_240_module_data_in[4] ;
 wire \sw_240_module_data_in[5] ;
 wire \sw_240_module_data_in[6] ;
 wire \sw_240_module_data_in[7] ;
 wire \sw_240_module_data_out[0] ;
 wire \sw_240_module_data_out[1] ;
 wire \sw_240_module_data_out[2] ;
 wire \sw_240_module_data_out[3] ;
 wire \sw_240_module_data_out[4] ;
 wire \sw_240_module_data_out[5] ;
 wire \sw_240_module_data_out[6] ;
 wire \sw_240_module_data_out[7] ;
 wire sw_240_scan_out;
 wire sw_241_clk_out;
 wire sw_241_data_out;
 wire sw_241_latch_out;
 wire \sw_241_module_data_in[0] ;
 wire \sw_241_module_data_in[1] ;
 wire \sw_241_module_data_in[2] ;
 wire \sw_241_module_data_in[3] ;
 wire \sw_241_module_data_in[4] ;
 wire \sw_241_module_data_in[5] ;
 wire \sw_241_module_data_in[6] ;
 wire \sw_241_module_data_in[7] ;
 wire \sw_241_module_data_out[0] ;
 wire \sw_241_module_data_out[1] ;
 wire \sw_241_module_data_out[2] ;
 wire \sw_241_module_data_out[3] ;
 wire \sw_241_module_data_out[4] ;
 wire \sw_241_module_data_out[5] ;
 wire \sw_241_module_data_out[6] ;
 wire \sw_241_module_data_out[7] ;
 wire sw_241_scan_out;
 wire sw_242_clk_out;
 wire sw_242_data_out;
 wire sw_242_latch_out;
 wire \sw_242_module_data_in[0] ;
 wire \sw_242_module_data_in[1] ;
 wire \sw_242_module_data_in[2] ;
 wire \sw_242_module_data_in[3] ;
 wire \sw_242_module_data_in[4] ;
 wire \sw_242_module_data_in[5] ;
 wire \sw_242_module_data_in[6] ;
 wire \sw_242_module_data_in[7] ;
 wire \sw_242_module_data_out[0] ;
 wire \sw_242_module_data_out[1] ;
 wire \sw_242_module_data_out[2] ;
 wire \sw_242_module_data_out[3] ;
 wire \sw_242_module_data_out[4] ;
 wire \sw_242_module_data_out[5] ;
 wire \sw_242_module_data_out[6] ;
 wire \sw_242_module_data_out[7] ;
 wire sw_242_scan_out;
 wire sw_243_clk_out;
 wire sw_243_data_out;
 wire sw_243_latch_out;
 wire \sw_243_module_data_in[0] ;
 wire \sw_243_module_data_in[1] ;
 wire \sw_243_module_data_in[2] ;
 wire \sw_243_module_data_in[3] ;
 wire \sw_243_module_data_in[4] ;
 wire \sw_243_module_data_in[5] ;
 wire \sw_243_module_data_in[6] ;
 wire \sw_243_module_data_in[7] ;
 wire \sw_243_module_data_out[0] ;
 wire \sw_243_module_data_out[1] ;
 wire \sw_243_module_data_out[2] ;
 wire \sw_243_module_data_out[3] ;
 wire \sw_243_module_data_out[4] ;
 wire \sw_243_module_data_out[5] ;
 wire \sw_243_module_data_out[6] ;
 wire \sw_243_module_data_out[7] ;
 wire sw_243_scan_out;
 wire sw_244_clk_out;
 wire sw_244_data_out;
 wire sw_244_latch_out;
 wire \sw_244_module_data_in[0] ;
 wire \sw_244_module_data_in[1] ;
 wire \sw_244_module_data_in[2] ;
 wire \sw_244_module_data_in[3] ;
 wire \sw_244_module_data_in[4] ;
 wire \sw_244_module_data_in[5] ;
 wire \sw_244_module_data_in[6] ;
 wire \sw_244_module_data_in[7] ;
 wire \sw_244_module_data_out[0] ;
 wire \sw_244_module_data_out[1] ;
 wire \sw_244_module_data_out[2] ;
 wire \sw_244_module_data_out[3] ;
 wire \sw_244_module_data_out[4] ;
 wire \sw_244_module_data_out[5] ;
 wire \sw_244_module_data_out[6] ;
 wire \sw_244_module_data_out[7] ;
 wire sw_244_scan_out;
 wire sw_245_clk_out;
 wire sw_245_data_out;
 wire sw_245_latch_out;
 wire \sw_245_module_data_in[0] ;
 wire \sw_245_module_data_in[1] ;
 wire \sw_245_module_data_in[2] ;
 wire \sw_245_module_data_in[3] ;
 wire \sw_245_module_data_in[4] ;
 wire \sw_245_module_data_in[5] ;
 wire \sw_245_module_data_in[6] ;
 wire \sw_245_module_data_in[7] ;
 wire \sw_245_module_data_out[0] ;
 wire \sw_245_module_data_out[1] ;
 wire \sw_245_module_data_out[2] ;
 wire \sw_245_module_data_out[3] ;
 wire \sw_245_module_data_out[4] ;
 wire \sw_245_module_data_out[5] ;
 wire \sw_245_module_data_out[6] ;
 wire \sw_245_module_data_out[7] ;
 wire sw_245_scan_out;
 wire sw_246_clk_out;
 wire sw_246_data_out;
 wire sw_246_latch_out;
 wire \sw_246_module_data_in[0] ;
 wire \sw_246_module_data_in[1] ;
 wire \sw_246_module_data_in[2] ;
 wire \sw_246_module_data_in[3] ;
 wire \sw_246_module_data_in[4] ;
 wire \sw_246_module_data_in[5] ;
 wire \sw_246_module_data_in[6] ;
 wire \sw_246_module_data_in[7] ;
 wire \sw_246_module_data_out[0] ;
 wire \sw_246_module_data_out[1] ;
 wire \sw_246_module_data_out[2] ;
 wire \sw_246_module_data_out[3] ;
 wire \sw_246_module_data_out[4] ;
 wire \sw_246_module_data_out[5] ;
 wire \sw_246_module_data_out[6] ;
 wire \sw_246_module_data_out[7] ;
 wire sw_246_scan_out;
 wire sw_247_clk_out;
 wire sw_247_data_out;
 wire sw_247_latch_out;
 wire \sw_247_module_data_in[0] ;
 wire \sw_247_module_data_in[1] ;
 wire \sw_247_module_data_in[2] ;
 wire \sw_247_module_data_in[3] ;
 wire \sw_247_module_data_in[4] ;
 wire \sw_247_module_data_in[5] ;
 wire \sw_247_module_data_in[6] ;
 wire \sw_247_module_data_in[7] ;
 wire \sw_247_module_data_out[0] ;
 wire \sw_247_module_data_out[1] ;
 wire \sw_247_module_data_out[2] ;
 wire \sw_247_module_data_out[3] ;
 wire \sw_247_module_data_out[4] ;
 wire \sw_247_module_data_out[5] ;
 wire \sw_247_module_data_out[6] ;
 wire \sw_247_module_data_out[7] ;
 wire sw_247_scan_out;
 wire sw_248_clk_out;
 wire sw_248_data_out;
 wire sw_248_latch_out;
 wire \sw_248_module_data_in[0] ;
 wire \sw_248_module_data_in[1] ;
 wire \sw_248_module_data_in[2] ;
 wire \sw_248_module_data_in[3] ;
 wire \sw_248_module_data_in[4] ;
 wire \sw_248_module_data_in[5] ;
 wire \sw_248_module_data_in[6] ;
 wire \sw_248_module_data_in[7] ;
 wire \sw_248_module_data_out[0] ;
 wire \sw_248_module_data_out[1] ;
 wire \sw_248_module_data_out[2] ;
 wire \sw_248_module_data_out[3] ;
 wire \sw_248_module_data_out[4] ;
 wire \sw_248_module_data_out[5] ;
 wire \sw_248_module_data_out[6] ;
 wire \sw_248_module_data_out[7] ;
 wire sw_248_scan_out;
 wire sw_249_latch_out;
 wire \sw_249_module_data_in[0] ;
 wire \sw_249_module_data_in[1] ;
 wire \sw_249_module_data_in[2] ;
 wire \sw_249_module_data_in[3] ;
 wire \sw_249_module_data_in[4] ;
 wire \sw_249_module_data_in[5] ;
 wire \sw_249_module_data_in[6] ;
 wire \sw_249_module_data_in[7] ;
 wire \sw_249_module_data_out[0] ;
 wire \sw_249_module_data_out[1] ;
 wire \sw_249_module_data_out[2] ;
 wire \sw_249_module_data_out[3] ;
 wire \sw_249_module_data_out[4] ;
 wire \sw_249_module_data_out[5] ;
 wire \sw_249_module_data_out[6] ;
 wire \sw_249_module_data_out[7] ;
 wire sw_249_scan_out;

 AidanMedcalf_pid_controller AidanMedcalf_pid_controller_076 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_076_module_data_in[7] ,
    \sw_076_module_data_in[6] ,
    \sw_076_module_data_in[5] ,
    \sw_076_module_data_in[4] ,
    \sw_076_module_data_in[3] ,
    \sw_076_module_data_in[2] ,
    \sw_076_module_data_in[1] ,
    \sw_076_module_data_in[0] }),
    .io_out({\sw_076_module_data_out[7] ,
    \sw_076_module_data_out[6] ,
    \sw_076_module_data_out[5] ,
    \sw_076_module_data_out[4] ,
    \sw_076_module_data_out[3] ,
    \sw_076_module_data_out[2] ,
    \sw_076_module_data_out[1] ,
    \sw_076_module_data_out[0] }));
 Asma_Mohsin_conv_enc_core Asma_Mohsin_conv_enc_core_118 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_118_module_data_in[7] ,
    \sw_118_module_data_in[6] ,
    \sw_118_module_data_in[5] ,
    \sw_118_module_data_in[4] ,
    \sw_118_module_data_in[3] ,
    \sw_118_module_data_in[2] ,
    \sw_118_module_data_in[1] ,
    \sw_118_module_data_in[0] }),
    .io_out({\sw_118_module_data_out[7] ,
    \sw_118_module_data_out[6] ,
    \sw_118_module_data_out[5] ,
    \sw_118_module_data_out[4] ,
    \sw_118_module_data_out[3] ,
    \sw_118_module_data_out[2] ,
    \sw_118_module_data_out[1] ,
    \sw_118_module_data_out[0] }));
 adamgreig_tt02_adc_dac adamgreig_tt02_adc_dac_100 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_100_module_data_in[7] ,
    \sw_100_module_data_in[6] ,
    \sw_100_module_data_in[5] ,
    \sw_100_module_data_in[4] ,
    \sw_100_module_data_in[3] ,
    \sw_100_module_data_in[2] ,
    \sw_100_module_data_in[1] ,
    \sw_100_module_data_in[0] }),
    .io_out({\sw_100_module_data_out[7] ,
    \sw_100_module_data_out[6] ,
    \sw_100_module_data_out[5] ,
    \sw_100_module_data_out[4] ,
    \sw_100_module_data_out[3] ,
    \sw_100_module_data_out[2] ,
    \sw_100_module_data_out[1] ,
    \sw_100_module_data_out[0] }));
 adamgreig_tt02_gps_ca_prn adamgreig_tt02_gps_ca_prn_099 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_099_module_data_in[7] ,
    \sw_099_module_data_in[6] ,
    \sw_099_module_data_in[5] ,
    \sw_099_module_data_in[4] ,
    \sw_099_module_data_in[3] ,
    \sw_099_module_data_in[2] ,
    \sw_099_module_data_in[1] ,
    \sw_099_module_data_in[0] }),
    .io_out({\sw_099_module_data_out[7] ,
    \sw_099_module_data_out[6] ,
    \sw_099_module_data_out[5] ,
    \sw_099_module_data_out[4] ,
    \sw_099_module_data_out[3] ,
    \sw_099_module_data_out[2] ,
    \sw_099_module_data_out[1] ,
    \sw_099_module_data_out[0] }));
 afoote_w5s8_tt02_top afoote_w5s8_tt02_top_125 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_125_module_data_in[7] ,
    \sw_125_module_data_in[6] ,
    \sw_125_module_data_in[5] ,
    \sw_125_module_data_in[4] ,
    \sw_125_module_data_in[3] ,
    \sw_125_module_data_in[2] ,
    \sw_125_module_data_in[1] ,
    \sw_125_module_data_in[0] }),
    .io_out({\sw_125_module_data_out[7] ,
    \sw_125_module_data_out[6] ,
    \sw_125_module_data_out[5] ,
    \sw_125_module_data_out[4] ,
    \sw_125_module_data_out[3] ,
    \sw_125_module_data_out[2] ,
    \sw_125_module_data_out[1] ,
    \sw_125_module_data_out[0] }));
 aidan_McCoy aidan_McCoy_008 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_008_module_data_in[7] ,
    \sw_008_module_data_in[6] ,
    \sw_008_module_data_in[5] ,
    \sw_008_module_data_in[4] ,
    \sw_008_module_data_in[3] ,
    \sw_008_module_data_in[2] ,
    \sw_008_module_data_in[1] ,
    \sw_008_module_data_in[0] }),
    .io_out({\sw_008_module_data_out[7] ,
    \sw_008_module_data_out[6] ,
    \sw_008_module_data_out[5] ,
    \sw_008_module_data_out[4] ,
    \sw_008_module_data_out[3] ,
    \sw_008_module_data_out[2] ,
    \sw_008_module_data_out[1] ,
    \sw_008_module_data_out[0] }));
 alu_top alu_top_007 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_007_module_data_in[7] ,
    \sw_007_module_data_in[6] ,
    \sw_007_module_data_in[5] ,
    \sw_007_module_data_in[4] ,
    \sw_007_module_data_in[3] ,
    \sw_007_module_data_in[2] ,
    \sw_007_module_data_in[1] ,
    \sw_007_module_data_in[0] }),
    .io_out({\sw_007_module_data_out[7] ,
    \sw_007_module_data_out[6] ,
    \sw_007_module_data_out[5] ,
    \sw_007_module_data_out[4] ,
    \sw_007_module_data_out[3] ,
    \sw_007_module_data_out[2] ,
    \sw_007_module_data_out[1] ,
    \sw_007_module_data_out[0] }));
 aramsey118_freq_counter aramsey118_freq_counter_088 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_088_module_data_in[7] ,
    \sw_088_module_data_in[6] ,
    \sw_088_module_data_in[5] ,
    \sw_088_module_data_in[4] ,
    \sw_088_module_data_in[3] ,
    \sw_088_module_data_in[2] ,
    \sw_088_module_data_in[1] ,
    \sw_088_module_data_in[0] }),
    .io_out({\sw_088_module_data_out[7] ,
    \sw_088_module_data_out[6] ,
    \sw_088_module_data_out[5] ,
    \sw_088_module_data_out[4] ,
    \sw_088_module_data_out[3] ,
    \sw_088_module_data_out[2] ,
    \sw_088_module_data_out[1] ,
    \sw_088_module_data_out[0] }));
 asic_multiplier_wrapper asic_multiplier_wrapper_023 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_023_module_data_in[7] ,
    \sw_023_module_data_in[6] ,
    \sw_023_module_data_in[5] ,
    \sw_023_module_data_in[4] ,
    \sw_023_module_data_in[3] ,
    \sw_023_module_data_in[2] ,
    \sw_023_module_data_in[1] ,
    \sw_023_module_data_in[0] }),
    .io_out({\sw_023_module_data_out[7] ,
    \sw_023_module_data_out[6] ,
    \sw_023_module_data_out[5] ,
    \sw_023_module_data_out[4] ,
    \sw_023_module_data_out[3] ,
    \sw_023_module_data_out[2] ,
    \sw_023_module_data_out[1] ,
    \sw_023_module_data_out[0] }));
 asinghani_beepboop asinghani_beepboop_151 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_151_module_data_in[7] ,
    \sw_151_module_data_in[6] ,
    \sw_151_module_data_in[5] ,
    \sw_151_module_data_in[4] ,
    \sw_151_module_data_in[3] ,
    \sw_151_module_data_in[2] ,
    \sw_151_module_data_in[1] ,
    \sw_151_module_data_in[0] }),
    .io_out({\sw_151_module_data_out[7] ,
    \sw_151_module_data_out[6] ,
    \sw_151_module_data_out[5] ,
    \sw_151_module_data_out[4] ,
    \sw_151_module_data_out[3] ,
    \sw_151_module_data_out[2] ,
    \sw_151_module_data_out[1] ,
    \sw_151_module_data_out[0] }));
 azdle_binary_clock azdle_binary_clock_009 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_009_module_data_in[7] ,
    \sw_009_module_data_in[6] ,
    \sw_009_module_data_in[5] ,
    \sw_009_module_data_in[4] ,
    \sw_009_module_data_in[3] ,
    \sw_009_module_data_in[2] ,
    \sw_009_module_data_in[1] ,
    \sw_009_module_data_in[0] }),
    .io_out({\sw_009_module_data_out[7] ,
    \sw_009_module_data_out[6] ,
    \sw_009_module_data_out[5] ,
    \sw_009_module_data_out[4] ,
    \sw_009_module_data_out[3] ,
    \sw_009_module_data_out[2] ,
    \sw_009_module_data_out[1] ,
    \sw_009_module_data_out[0] }));
 browndeer_rv8u browndeer_rv8u_107 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_107_module_data_in[7] ,
    \sw_107_module_data_in[6] ,
    \sw_107_module_data_in[5] ,
    \sw_107_module_data_in[4] ,
    \sw_107_module_data_in[3] ,
    \sw_107_module_data_in[2] ,
    \sw_107_module_data_in[1] ,
    \sw_107_module_data_in[0] }),
    .io_out({\sw_107_module_data_out[7] ,
    \sw_107_module_data_out[6] ,
    \sw_107_module_data_out[5] ,
    \sw_107_module_data_out[4] ,
    \sw_107_module_data_out[3] ,
    \sw_107_module_data_out[2] ,
    \sw_107_module_data_out[1] ,
    \sw_107_module_data_out[0] }));
 cchan_fp8_multiplier cchan_fp8_multiplier_060 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_060_module_data_in[7] ,
    \sw_060_module_data_in[6] ,
    \sw_060_module_data_in[5] ,
    \sw_060_module_data_in[4] ,
    \sw_060_module_data_in[3] ,
    \sw_060_module_data_in[2] ,
    \sw_060_module_data_in[1] ,
    \sw_060_module_data_in[0] }),
    .io_out({\sw_060_module_data_out[7] ,
    \sw_060_module_data_out[6] ,
    \sw_060_module_data_out[5] ,
    \sw_060_module_data_out[4] ,
    \sw_060_module_data_out[3] ,
    \sw_060_module_data_out[2] ,
    \sw_060_module_data_out[1] ,
    \sw_060_module_data_out[0] }));
 chase_the_beat chase_the_beat_020 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_020_module_data_in[7] ,
    \sw_020_module_data_in[6] ,
    \sw_020_module_data_in[5] ,
    \sw_020_module_data_in[4] ,
    \sw_020_module_data_in[3] ,
    \sw_020_module_data_in[2] ,
    \sw_020_module_data_in[1] ,
    \sw_020_module_data_in[0] }),
    .io_out({\sw_020_module_data_out[7] ,
    \sw_020_module_data_out[6] ,
    \sw_020_module_data_out[5] ,
    \sw_020_module_data_out[4] ,
    \sw_020_module_data_out[3] ,
    \sw_020_module_data_out[2] ,
    \sw_020_module_data_out[1] ,
    \sw_020_module_data_out[0] }));
 chrisruk_matrix chrisruk_matrix_003 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_003_module_data_in[7] ,
    \sw_003_module_data_in[6] ,
    \sw_003_module_data_in[5] ,
    \sw_003_module_data_in[4] ,
    \sw_003_module_data_in[3] ,
    \sw_003_module_data_in[2] ,
    \sw_003_module_data_in[1] ,
    \sw_003_module_data_in[0] }),
    .io_out({\sw_003_module_data_out[7] ,
    \sw_003_module_data_out[6] ,
    \sw_003_module_data_out[5] ,
    \sw_003_module_data_out[4] ,
    \sw_003_module_data_out[3] ,
    \sw_003_module_data_out[2] ,
    \sw_003_module_data_out[1] ,
    \sw_003_module_data_out[0] }));
 cpldcpu_MCPU5plus cpldcpu_MCPU5plus_078 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_078_module_data_in[7] ,
    \sw_078_module_data_in[6] ,
    \sw_078_module_data_in[5] ,
    \sw_078_module_data_in[4] ,
    \sw_078_module_data_in[3] ,
    \sw_078_module_data_in[2] ,
    \sw_078_module_data_in[1] ,
    \sw_078_module_data_in[0] }),
    .io_out({\sw_078_module_data_out[7] ,
    \sw_078_module_data_out[6] ,
    \sw_078_module_data_out[5] ,
    \sw_078_module_data_out[4] ,
    \sw_078_module_data_out[3] ,
    \sw_078_module_data_out[2] ,
    \sw_078_module_data_out[1] ,
    \sw_078_module_data_out[0] }));
 cpldcpu_TrainLED2top cpldcpu_TrainLED2top_077 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_077_module_data_in[7] ,
    \sw_077_module_data_in[6] ,
    \sw_077_module_data_in[5] ,
    \sw_077_module_data_in[4] ,
    \sw_077_module_data_in[3] ,
    \sw_077_module_data_in[2] ,
    \sw_077_module_data_in[1] ,
    \sw_077_module_data_in[0] }),
    .io_out({\sw_077_module_data_out[7] ,
    \sw_077_module_data_out[6] ,
    \sw_077_module_data_out[5] ,
    \sw_077_module_data_out[4] ,
    \sw_077_module_data_out[3] ,
    \sw_077_module_data_out[2] ,
    \sw_077_module_data_out[1] ,
    \sw_077_module_data_out[0] }));
 davidsiaw_stackcalc davidsiaw_stackcalc_080 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_080_module_data_in[7] ,
    \sw_080_module_data_in[6] ,
    \sw_080_module_data_in[5] ,
    \sw_080_module_data_in[4] ,
    \sw_080_module_data_in[3] ,
    \sw_080_module_data_in[2] ,
    \sw_080_module_data_in[1] ,
    \sw_080_module_data_in[0] }),
    .io_out({\sw_080_module_data_out[7] ,
    \sw_080_module_data_out[6] ,
    \sw_080_module_data_out[5] ,
    \sw_080_module_data_out[4] ,
    \sw_080_module_data_out[3] ,
    \sw_080_module_data_out[2] ,
    \sw_080_module_data_out[1] ,
    \sw_080_module_data_out[0] }));
 ericsmi_speed_test ericsmi_speed_test_075 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_075_module_data_in[7] ,
    \sw_075_module_data_in[6] ,
    \sw_075_module_data_in[5] ,
    \sw_075_module_data_in[4] ,
    \sw_075_module_data_in[3] ,
    \sw_075_module_data_in[2] ,
    \sw_075_module_data_in[1] ,
    \sw_075_module_data_in[0] }),
    .io_out({\sw_075_module_data_out[7] ,
    \sw_075_module_data_out[6] ,
    \sw_075_module_data_out[5] ,
    \sw_075_module_data_out[4] ,
    \sw_075_module_data_out[3] ,
    \sw_075_module_data_out[2] ,
    \sw_075_module_data_out[1] ,
    \sw_075_module_data_out[0] }));
 femto_top femto_top_143 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_143_module_data_in[7] ,
    \sw_143_module_data_in[6] ,
    \sw_143_module_data_in[5] ,
    \sw_143_module_data_in[4] ,
    \sw_143_module_data_in[3] ,
    \sw_143_module_data_in[2] ,
    \sw_143_module_data_in[1] ,
    \sw_143_module_data_in[0] }),
    .io_out({\sw_143_module_data_out[7] ,
    \sw_143_module_data_out[6] ,
    \sw_143_module_data_out[5] ,
    \sw_143_module_data_out[4] ,
    \sw_143_module_data_out[3] ,
    \sw_143_module_data_out[2] ,
    \sw_143_module_data_out[1] ,
    \sw_143_module_data_out[0] }));
 flygoat_tt02_play_tune flygoat_tt02_play_tune_054 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_054_module_data_in[7] ,
    \sw_054_module_data_in[6] ,
    \sw_054_module_data_in[5] ,
    \sw_054_module_data_in[4] ,
    \sw_054_module_data_in[3] ,
    \sw_054_module_data_in[2] ,
    \sw_054_module_data_in[1] ,
    \sw_054_module_data_in[0] }),
    .io_out({\sw_054_module_data_out[7] ,
    \sw_054_module_data_out[6] ,
    \sw_054_module_data_out[5] ,
    \sw_054_module_data_out[4] ,
    \sw_054_module_data_out[3] ,
    \sw_054_module_data_out[2] ,
    \sw_054_module_data_out[1] ,
    \sw_054_module_data_out[0] }));
 fraserbc_simon fraserbc_simon_001 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_001_module_data_in[7] ,
    \sw_001_module_data_in[6] ,
    \sw_001_module_data_in[5] ,
    \sw_001_module_data_in[4] ,
    \sw_001_module_data_in[3] ,
    \sw_001_module_data_in[2] ,
    \sw_001_module_data_in[1] ,
    \sw_001_module_data_in[0] }),
    .io_out({\sw_001_module_data_out[7] ,
    \sw_001_module_data_out[6] ,
    \sw_001_module_data_out[5] ,
    \sw_001_module_data_out[4] ,
    \sw_001_module_data_out[3] ,
    \sw_001_module_data_out[2] ,
    \sw_001_module_data_out[1] ,
    \sw_001_module_data_out[0] }));
 frog frog_114 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_114_module_data_in[7] ,
    \sw_114_module_data_in[6] ,
    \sw_114_module_data_in[5] ,
    \sw_114_module_data_in[4] ,
    \sw_114_module_data_in[3] ,
    \sw_114_module_data_in[2] ,
    \sw_114_module_data_in[1] ,
    \sw_114_module_data_in[0] }),
    .io_out({\sw_114_module_data_out[7] ,
    \sw_114_module_data_out[6] ,
    \sw_114_module_data_out[5] ,
    \sw_114_module_data_out[4] ,
    \sw_114_module_data_out[3] ,
    \sw_114_module_data_out[2] ,
    \sw_114_module_data_out[1] ,
    \sw_114_module_data_out[0] }));
 gatecat_fpga_top gatecat_fpga_top_090 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_090_module_data_in[7] ,
    \sw_090_module_data_in[6] ,
    \sw_090_module_data_in[5] ,
    \sw_090_module_data_in[4] ,
    \sw_090_module_data_in[3] ,
    \sw_090_module_data_in[2] ,
    \sw_090_module_data_in[1] ,
    \sw_090_module_data_in[0] }),
    .io_out({\sw_090_module_data_out[7] ,
    \sw_090_module_data_out[6] ,
    \sw_090_module_data_out[5] ,
    \sw_090_module_data_out[4] ,
    \sw_090_module_data_out[3] ,
    \sw_090_module_data_out[2] ,
    \sw_090_module_data_out[1] ,
    \sw_090_module_data_out[0] }));
 github_com_proppy_tt02_xls_counter github_com_proppy_tt02_xls_counter_051 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_051_module_data_in[7] ,
    \sw_051_module_data_in[6] ,
    \sw_051_module_data_in[5] ,
    \sw_051_module_data_in[4] ,
    \sw_051_module_data_in[3] ,
    \sw_051_module_data_in[2] ,
    \sw_051_module_data_in[1] ,
    \sw_051_module_data_in[0] }),
    .io_out({\sw_051_module_data_out[7] ,
    \sw_051_module_data_out[6] ,
    \sw_051_module_data_out[5] ,
    \sw_051_module_data_out[4] ,
    \sw_051_module_data_out[3] ,
    \sw_051_module_data_out[2] ,
    \sw_051_module_data_out[1] ,
    \sw_051_module_data_out[0] }));
 github_com_proppy_tt02_xls_popcount github_com_proppy_tt02_xls_popcount_042 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_042_module_data_in[7] ,
    \sw_042_module_data_in[6] ,
    \sw_042_module_data_in[5] ,
    \sw_042_module_data_in[4] ,
    \sw_042_module_data_in[3] ,
    \sw_042_module_data_in[2] ,
    \sw_042_module_data_in[1] ,
    \sw_042_module_data_in[0] }),
    .io_out({\sw_042_module_data_out[7] ,
    \sw_042_module_data_out[6] ,
    \sw_042_module_data_out[5] ,
    \sw_042_module_data_out[4] ,
    \sw_042_module_data_out[3] ,
    \sw_042_module_data_out[2] ,
    \sw_042_module_data_out[1] ,
    \sw_042_module_data_out[0] }));
 gregdavill_clock_top gregdavill_clock_top_127 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_127_module_data_in[7] ,
    \sw_127_module_data_in[6] ,
    \sw_127_module_data_in[5] ,
    \sw_127_module_data_in[4] ,
    \sw_127_module_data_in[3] ,
    \sw_127_module_data_in[2] ,
    \sw_127_module_data_in[1] ,
    \sw_127_module_data_in[0] }),
    .io_out({\sw_127_module_data_out[7] ,
    \sw_127_module_data_out[6] ,
    \sw_127_module_data_out[5] ,
    \sw_127_module_data_out[4] ,
    \sw_127_module_data_out[3] ,
    \sw_127_module_data_out[2] ,
    \sw_127_module_data_out[1] ,
    \sw_127_module_data_out[0] }));
 gregdavill_serv_top gregdavill_serv_top_128 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_128_module_data_in[7] ,
    \sw_128_module_data_in[6] ,
    \sw_128_module_data_in[5] ,
    \sw_128_module_data_in[4] ,
    \sw_128_module_data_in[3] ,
    \sw_128_module_data_in[2] ,
    \sw_128_module_data_in[1] ,
    \sw_128_module_data_in[0] }),
    .io_out({\sw_128_module_data_out[7] ,
    \sw_128_module_data_out[6] ,
    \sw_128_module_data_out[5] ,
    \sw_128_module_data_out[4] ,
    \sw_128_module_data_out[3] ,
    \sw_128_module_data_out[2] ,
    \sw_128_module_data_out[1] ,
    \sw_128_module_data_out[0] }));
 hex_sr hex_sr_074 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_074_module_data_in[7] ,
    \sw_074_module_data_in[6] ,
    \sw_074_module_data_in[5] ,
    \sw_074_module_data_in[4] ,
    \sw_074_module_data_in[3] ,
    \sw_074_module_data_in[2] ,
    \sw_074_module_data_in[1] ,
    \sw_074_module_data_in[0] }),
    .io_out({\sw_074_module_data_out[7] ,
    \sw_074_module_data_out[6] ,
    \sw_074_module_data_out[5] ,
    \sw_074_module_data_out[4] ,
    \sw_074_module_data_out[3] ,
    \sw_074_module_data_out[2] ,
    \sw_074_module_data_out[1] ,
    \sw_074_module_data_out[0] }));
 jar_pi jar_pi_036 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_036_module_data_in[7] ,
    \sw_036_module_data_in[6] ,
    \sw_036_module_data_in[5] ,
    \sw_036_module_data_in[4] ,
    \sw_036_module_data_in[3] ,
    \sw_036_module_data_in[2] ,
    \sw_036_module_data_in[1] ,
    \sw_036_module_data_in[0] }),
    .io_out({\sw_036_module_data_out[7] ,
    \sw_036_module_data_out[6] ,
    \sw_036_module_data_out[5] ,
    \sw_036_module_data_out[4] ,
    \sw_036_module_data_out[3] ,
    \sw_036_module_data_out[2] ,
    \sw_036_module_data_out[1] ,
    \sw_036_module_data_out[0] }));
 jar_sram_top jar_sram_top_011 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_011_module_data_in[7] ,
    \sw_011_module_data_in[6] ,
    \sw_011_module_data_in[5] ,
    \sw_011_module_data_in[4] ,
    \sw_011_module_data_in[3] ,
    \sw_011_module_data_in[2] ,
    \sw_011_module_data_in[1] ,
    \sw_011_module_data_in[0] }),
    .io_out({\sw_011_module_data_out[7] ,
    \sw_011_module_data_out[6] ,
    \sw_011_module_data_out[5] ,
    \sw_011_module_data_out[4] ,
    \sw_011_module_data_out[3] ,
    \sw_011_module_data_out[2] ,
    \sw_011_module_data_out[1] ,
    \sw_011_module_data_out[0] }));
 jglim_7seg jglim_7seg_101 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_101_module_data_in[7] ,
    \sw_101_module_data_in[6] ,
    \sw_101_module_data_in[5] ,
    \sw_101_module_data_in[4] ,
    \sw_101_module_data_in[3] ,
    \sw_101_module_data_in[2] ,
    \sw_101_module_data_in[1] ,
    \sw_101_module_data_in[0] }),
    .io_out({\sw_101_module_data_out[7] ,
    \sw_101_module_data_out[6] ,
    \sw_101_module_data_out[5] ,
    \sw_101_module_data_out[4] ,
    \sw_101_module_data_out[3] ,
    \sw_101_module_data_out[2] ,
    \sw_101_module_data_out[1] ,
    \sw_101_module_data_out[0] }));
 jleightcap_top jleightcap_top_055 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_055_module_data_in[7] ,
    \sw_055_module_data_in[6] ,
    \sw_055_module_data_in[5] ,
    \sw_055_module_data_in[4] ,
    \sw_055_module_data_in[3] ,
    \sw_055_module_data_in[2] ,
    \sw_055_module_data_in[1] ,
    \sw_055_module_data_in[0] }),
    .io_out({\sw_055_module_data_out[7] ,
    \sw_055_module_data_out[6] ,
    \sw_055_module_data_out[5] ,
    \sw_055_module_data_out[4] ,
    \sw_055_module_data_out[3] ,
    \sw_055_module_data_out[2] ,
    \sw_055_module_data_out[1] ,
    \sw_055_module_data_out[0] }));
 jonpaolo02_async_fifo jonpaolo02_async_fifo_150 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_150_module_data_in[7] ,
    \sw_150_module_data_in[6] ,
    \sw_150_module_data_in[5] ,
    \sw_150_module_data_in[4] ,
    \sw_150_module_data_in[3] ,
    \sw_150_module_data_in[2] ,
    \sw_150_module_data_in[1] ,
    \sw_150_module_data_in[0] }),
    .io_out({\sw_150_module_data_out[7] ,
    \sw_150_module_data_out[6] ,
    \sw_150_module_data_out[5] ,
    \sw_150_module_data_out[4] ,
    \sw_150_module_data_out[3] ,
    \sw_150_module_data_out[2] ,
    \sw_150_module_data_out[1] ,
    \sw_150_module_data_out[0] }));
 klei22_ra klei22_ra_124 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_124_module_data_in[7] ,
    \sw_124_module_data_in[6] ,
    \sw_124_module_data_in[5] ,
    \sw_124_module_data_in[4] ,
    \sw_124_module_data_in[3] ,
    \sw_124_module_data_in[2] ,
    \sw_124_module_data_in[1] ,
    \sw_124_module_data_in[0] }),
    .io_out({\sw_124_module_data_out[7] ,
    \sw_124_module_data_out[6] ,
    \sw_124_module_data_out[5] ,
    \sw_124_module_data_out[4] ,
    \sw_124_module_data_out[3] ,
    \sw_124_module_data_out[2] ,
    \sw_124_module_data_out[1] ,
    \sw_124_module_data_out[0] }));
 krasin_3_bit_8_channel_pwm_driver krasin_3_bit_8_channel_pwm_driver_058 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_058_module_data_in[7] ,
    \sw_058_module_data_in[6] ,
    \sw_058_module_data_in[5] ,
    \sw_058_module_data_in[4] ,
    \sw_058_module_data_in[3] ,
    \sw_058_module_data_in[2] ,
    \sw_058_module_data_in[1] ,
    \sw_058_module_data_in[0] }),
    .io_out({\sw_058_module_data_out[7] ,
    \sw_058_module_data_out[6] ,
    \sw_058_module_data_out[5] ,
    \sw_058_module_data_out[4] ,
    \sw_058_module_data_out[3] ,
    \sw_058_module_data_out[2] ,
    \sw_058_module_data_out[1] ,
    \sw_058_module_data_out[0] }));
 krasin_tt02_verilog_spi_7_channel_pwm_driver krasin_tt02_verilog_spi_7_channel_pwm_driver_073 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_073_module_data_in[7] ,
    \sw_073_module_data_in[6] ,
    \sw_073_module_data_in[5] ,
    \sw_073_module_data_in[4] ,
    \sw_073_module_data_in[3] ,
    \sw_073_module_data_in[2] ,
    \sw_073_module_data_in[1] ,
    \sw_073_module_data_in[0] }),
    .io_out({\sw_073_module_data_out[7] ,
    \sw_073_module_data_out[6] ,
    \sw_073_module_data_out[5] ,
    \sw_073_module_data_out[4] ,
    \sw_073_module_data_out[3] ,
    \sw_073_module_data_out[2] ,
    \sw_073_module_data_out[1] ,
    \sw_073_module_data_out[0] }));
 logisim_demo logisim_demo_144 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_144_module_data_in[7] ,
    \sw_144_module_data_in[6] ,
    \sw_144_module_data_in[5] ,
    \sw_144_module_data_in[4] ,
    \sw_144_module_data_in[3] ,
    \sw_144_module_data_in[2] ,
    \sw_144_module_data_in[1] ,
    \sw_144_module_data_in[0] }),
    .io_out({\sw_144_module_data_out[7] ,
    \sw_144_module_data_out[6] ,
    \sw_144_module_data_out[5] ,
    \sw_144_module_data_out[4] ,
    \sw_144_module_data_out[3] ,
    \sw_144_module_data_out[2] ,
    \sw_144_module_data_out[1] ,
    \sw_144_module_data_out[0] }));
 loxodes_sequencer loxodes_sequencer_004 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_004_module_data_in[7] ,
    \sw_004_module_data_in[6] ,
    \sw_004_module_data_in[5] ,
    \sw_004_module_data_in[4] ,
    \sw_004_module_data_in[3] ,
    \sw_004_module_data_in[2] ,
    \sw_004_module_data_in[1] ,
    \sw_004_module_data_in[0] }),
    .io_out({\sw_004_module_data_out[7] ,
    \sw_004_module_data_out[6] ,
    \sw_004_module_data_out[5] ,
    \sw_004_module_data_out[4] ,
    \sw_004_module_data_out[3] ,
    \sw_004_module_data_out[2] ,
    \sw_004_module_data_out[1] ,
    \sw_004_module_data_out[0] }));
 luthor2k_top_tto luthor2k_top_tto_116 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_116_module_data_in[7] ,
    \sw_116_module_data_in[6] ,
    \sw_116_module_data_in[5] ,
    \sw_116_module_data_in[4] ,
    \sw_116_module_data_in[3] ,
    \sw_116_module_data_in[2] ,
    \sw_116_module_data_in[1] ,
    \sw_116_module_data_in[0] }),
    .io_out({\sw_116_module_data_out[7] ,
    \sw_116_module_data_out[6] ,
    \sw_116_module_data_out[5] ,
    \sw_116_module_data_out[4] ,
    \sw_116_module_data_out[3] ,
    \sw_116_module_data_out[2] ,
    \sw_116_module_data_out[1] ,
    \sw_116_module_data_out[0] }));
 mbikovitsky_top mbikovitsky_top_033 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_033_module_data_in[7] ,
    \sw_033_module_data_in[6] ,
    \sw_033_module_data_in[5] ,
    \sw_033_module_data_in[4] ,
    \sw_033_module_data_in[3] ,
    \sw_033_module_data_in[2] ,
    \sw_033_module_data_in[1] ,
    \sw_033_module_data_in[0] }),
    .io_out({\sw_033_module_data_out[7] ,
    \sw_033_module_data_out[6] ,
    \sw_033_module_data_out[5] ,
    \sw_033_module_data_out[4] ,
    \sw_033_module_data_out[3] ,
    \sw_033_module_data_out[2] ,
    \sw_033_module_data_out[1] ,
    \sw_033_module_data_out[0] }));
 meriac_tt02_play_tune meriac_tt02_play_tune_045 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_045_module_data_in[7] ,
    \sw_045_module_data_in[6] ,
    \sw_045_module_data_in[5] ,
    \sw_045_module_data_in[4] ,
    \sw_045_module_data_in[3] ,
    \sw_045_module_data_in[2] ,
    \sw_045_module_data_in[1] ,
    \sw_045_module_data_in[0] }),
    .io_out({\sw_045_module_data_out[7] ,
    \sw_045_module_data_out[6] ,
    \sw_045_module_data_out[5] ,
    \sw_045_module_data_out[4] ,
    \sw_045_module_data_out[3] ,
    \sw_045_module_data_out[2] ,
    \sw_045_module_data_out[1] ,
    \sw_045_module_data_out[0] }));
 migcorre_pwm migcorre_pwm_005 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_005_module_data_in[7] ,
    \sw_005_module_data_in[6] ,
    \sw_005_module_data_in[5] ,
    \sw_005_module_data_in[4] ,
    \sw_005_module_data_in[3] ,
    \sw_005_module_data_in[2] ,
    \sw_005_module_data_in[1] ,
    \sw_005_module_data_in[0] }),
    .io_out({\sw_005_module_data_out[7] ,
    \sw_005_module_data_out[6] ,
    \sw_005_module_data_out[5] ,
    \sw_005_module_data_out[4] ,
    \sw_005_module_data_out[3] ,
    \sw_005_module_data_out[2] ,
    \sw_005_module_data_out[1] ,
    \sw_005_module_data_out[0] }));
 mm21_LEDMatrixTop mm21_LEDMatrixTop_026 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_026_module_data_in[7] ,
    \sw_026_module_data_in[6] ,
    \sw_026_module_data_in[5] ,
    \sw_026_module_data_in[4] ,
    \sw_026_module_data_in[3] ,
    \sw_026_module_data_in[2] ,
    \sw_026_module_data_in[1] ,
    \sw_026_module_data_in[0] }),
    .io_out({\sw_026_module_data_out[7] ,
    \sw_026_module_data_out[6] ,
    \sw_026_module_data_out[5] ,
    \sw_026_module_data_out[4] ,
    \sw_026_module_data_out[3] ,
    \sw_026_module_data_out[2] ,
    \sw_026_module_data_out[1] ,
    \sw_026_module_data_out[0] }));
 moonbase_cpu_4bit moonbase_cpu_4bit_079 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_079_module_data_in[7] ,
    \sw_079_module_data_in[6] ,
    \sw_079_module_data_in[5] ,
    \sw_079_module_data_in[4] ,
    \sw_079_module_data_in[3] ,
    \sw_079_module_data_in[2] ,
    \sw_079_module_data_in[1] ,
    \sw_079_module_data_in[0] }),
    .io_out({\sw_079_module_data_out[7] ,
    \sw_079_module_data_out[6] ,
    \sw_079_module_data_out[5] ,
    \sw_079_module_data_out[4] ,
    \sw_079_module_data_out[3] ,
    \sw_079_module_data_out[2] ,
    \sw_079_module_data_out[1] ,
    \sw_079_module_data_out[0] }));
 moonbase_cpu_8bit moonbase_cpu_8bit_085 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_085_module_data_in[7] ,
    \sw_085_module_data_in[6] ,
    \sw_085_module_data_in[5] ,
    \sw_085_module_data_in[4] ,
    \sw_085_module_data_in[3] ,
    \sw_085_module_data_in[2] ,
    \sw_085_module_data_in[1] ,
    \sw_085_module_data_in[0] }),
    .io_out({\sw_085_module_data_out[7] ,
    \sw_085_module_data_out[6] ,
    \sw_085_module_data_out[5] ,
    \sw_085_module_data_out[4] ,
    \sw_085_module_data_out[3] ,
    \sw_085_module_data_out[2] ,
    \sw_085_module_data_out[1] ,
    \sw_085_module_data_out[0] }));
 moyes0_top_module moyes0_top_module_039 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_039_module_data_in[7] ,
    \sw_039_module_data_in[6] ,
    \sw_039_module_data_in[5] ,
    \sw_039_module_data_in[4] ,
    \sw_039_module_data_in[3] ,
    \sw_039_module_data_in[2] ,
    \sw_039_module_data_in[1] ,
    \sw_039_module_data_in[0] }),
    .io_out({\sw_039_module_data_out[7] ,
    \sw_039_module_data_out[6] ,
    \sw_039_module_data_out[5] ,
    \sw_039_module_data_out[4] ,
    \sw_039_module_data_out[3] ,
    \sw_039_module_data_out[2] ,
    \sw_039_module_data_out[1] ,
    \sw_039_module_data_out[0] }));
 msaghir_top_level msaghir_top_level_135 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_135_module_data_in[7] ,
    \sw_135_module_data_in[6] ,
    \sw_135_module_data_in[5] ,
    \sw_135_module_data_in[4] ,
    \sw_135_module_data_in[3] ,
    \sw_135_module_data_in[2] ,
    \sw_135_module_data_in[1] ,
    \sw_135_module_data_in[0] }),
    .io_out({\sw_135_module_data_out[7] ,
    \sw_135_module_data_out[6] ,
    \sw_135_module_data_out[5] ,
    \sw_135_module_data_out[4] ,
    \sw_135_module_data_out[3] ,
    \sw_135_module_data_out[2] ,
    \sw_135_module_data_out[1] ,
    \sw_135_module_data_out[0] }));
 navray_top navray_top_071 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_071_module_data_in[7] ,
    \sw_071_module_data_in[6] ,
    \sw_071_module_data_in[5] ,
    \sw_071_module_data_in[4] ,
    \sw_071_module_data_in[3] ,
    \sw_071_module_data_in[2] ,
    \sw_071_module_data_in[1] ,
    \sw_071_module_data_in[0] }),
    .io_out({\sw_071_module_data_out[7] ,
    \sw_071_module_data_out[6] ,
    \sw_071_module_data_out[5] ,
    \sw_071_module_data_out[4] ,
    \sw_071_module_data_out[3] ,
    \sw_071_module_data_out[2] ,
    \sw_071_module_data_out[1] ,
    \sw_071_module_data_out[0] }));
 noahgaertner_cpu noahgaertner_cpu_152 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_152_module_data_in[7] ,
    \sw_152_module_data_in[6] ,
    \sw_152_module_data_in[5] ,
    \sw_152_module_data_in[4] ,
    \sw_152_module_data_in[3] ,
    \sw_152_module_data_in[2] ,
    \sw_152_module_data_in[1] ,
    \sw_152_module_data_in[0] }),
    .io_out({\sw_152_module_data_out[7] ,
    \sw_152_module_data_out[6] ,
    \sw_152_module_data_out[5] ,
    \sw_152_module_data_out[4] ,
    \sw_152_module_data_out[3] ,
    \sw_152_module_data_out[2] ,
    \sw_152_module_data_out[1] ,
    \sw_152_module_data_out[0] }));
 option22 option22_139 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_139_module_data_in[7] ,
    \sw_139_module_data_in[6] ,
    \sw_139_module_data_in[5] ,
    \sw_139_module_data_in[4] ,
    \sw_139_module_data_in[3] ,
    \sw_139_module_data_in[2] ,
    \sw_139_module_data_in[1] ,
    \sw_139_module_data_in[0] }),
    .io_out({\sw_139_module_data_out[7] ,
    \sw_139_module_data_out[6] ,
    \sw_139_module_data_out[5] ,
    \sw_139_module_data_out[4] ,
    \sw_139_module_data_out[3] ,
    \sw_139_module_data_out[2] ,
    \sw_139_module_data_out[1] ,
    \sw_139_module_data_out[0] }));
 option23 option23_138 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_138_module_data_in[7] ,
    \sw_138_module_data_in[6] ,
    \sw_138_module_data_in[5] ,
    \sw_138_module_data_in[4] ,
    \sw_138_module_data_in[3] ,
    \sw_138_module_data_in[2] ,
    \sw_138_module_data_in[1] ,
    \sw_138_module_data_in[0] }),
    .io_out({\sw_138_module_data_out[7] ,
    \sw_138_module_data_out[6] ,
    \sw_138_module_data_out[5] ,
    \sw_138_module_data_out[4] ,
    \sw_138_module_data_out[3] ,
    \sw_138_module_data_out[2] ,
    \sw_138_module_data_out[1] ,
    \sw_138_module_data_out[0] }));
 option23ser option23ser_137 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_137_module_data_in[7] ,
    \sw_137_module_data_in[6] ,
    \sw_137_module_data_in[5] ,
    \sw_137_module_data_in[4] ,
    \sw_137_module_data_in[3] ,
    \sw_137_module_data_in[2] ,
    \sw_137_module_data_in[1] ,
    \sw_137_module_data_in[0] }),
    .io_out({\sw_137_module_data_out[7] ,
    \sw_137_module_data_out[6] ,
    \sw_137_module_data_out[5] ,
    \sw_137_module_data_out[4] ,
    \sw_137_module_data_out[3] ,
    \sw_137_module_data_out[2] ,
    \sw_137_module_data_out[1] ,
    \sw_137_module_data_out[0] }));
 phasenoisepon_seven_segment_seconds phasenoisepon_seven_segment_seconds_046 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_046_module_data_in[7] ,
    \sw_046_module_data_in[6] ,
    \sw_046_module_data_in[5] ,
    \sw_046_module_data_in[4] ,
    \sw_046_module_data_in[3] ,
    \sw_046_module_data_in[2] ,
    \sw_046_module_data_in[1] ,
    \sw_046_module_data_in[0] }),
    .io_out({\sw_046_module_data_out[7] ,
    \sw_046_module_data_out[6] ,
    \sw_046_module_data_out[5] ,
    \sw_046_module_data_out[4] ,
    \sw_046_module_data_out[3] ,
    \sw_046_module_data_out[2] ,
    \sw_046_module_data_out[1] ,
    \sw_046_module_data_out[0] }));
 poisonninja_top poisonninja_top_147 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_147_module_data_in[7] ,
    \sw_147_module_data_in[6] ,
    \sw_147_module_data_in[5] ,
    \sw_147_module_data_in[4] ,
    \sw_147_module_data_in[3] ,
    \sw_147_module_data_in[2] ,
    \sw_147_module_data_in[1] ,
    \sw_147_module_data_in[0] }),
    .io_out({\sw_147_module_data_out[7] ,
    \sw_147_module_data_out[6] ,
    \sw_147_module_data_out[5] ,
    \sw_147_module_data_out[4] ,
    \sw_147_module_data_out[3] ,
    \sw_147_module_data_out[2] ,
    \sw_147_module_data_out[1] ,
    \sw_147_module_data_out[0] }));
 prog_melody_gen prog_melody_gen_109 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_109_module_data_in[7] ,
    \sw_109_module_data_in[6] ,
    \sw_109_module_data_in[5] ,
    \sw_109_module_data_in[4] ,
    \sw_109_module_data_in[3] ,
    \sw_109_module_data_in[2] ,
    \sw_109_module_data_in[1] ,
    \sw_109_module_data_in[0] }),
    .io_out({\sw_109_module_data_out[7] ,
    \sw_109_module_data_out[6] ,
    \sw_109_module_data_out[5] ,
    \sw_109_module_data_out[4] ,
    \sw_109_module_data_out[3] ,
    \sw_109_module_data_out[2] ,
    \sw_109_module_data_out[1] ,
    \sw_109_module_data_out[0] }));
 pwm_gen pwm_gen_068 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_068_module_data_in[7] ,
    \sw_068_module_data_in[6] ,
    \sw_068_module_data_in[5] ,
    \sw_068_module_data_in[4] ,
    \sw_068_module_data_in[3] ,
    \sw_068_module_data_in[2] ,
    \sw_068_module_data_in[1] ,
    \sw_068_module_data_in[0] }),
    .io_out({\sw_068_module_data_out[7] ,
    \sw_068_module_data_out[6] ,
    \sw_068_module_data_out[5] ,
    \sw_068_module_data_out[4] ,
    \sw_068_module_data_out[3] ,
    \sw_068_module_data_out[2] ,
    \sw_068_module_data_out[1] ,
    \sw_068_module_data_out[0] }));
 razhas_top_level razhas_top_level_164 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_164_module_data_in[7] ,
    \sw_164_module_data_in[6] ,
    \sw_164_module_data_in[5] ,
    \sw_164_module_data_in[4] ,
    \sw_164_module_data_in[3] ,
    \sw_164_module_data_in[2] ,
    \sw_164_module_data_in[1] ,
    \sw_164_module_data_in[0] }),
    .io_out({\sw_164_module_data_out[7] ,
    \sw_164_module_data_out[6] ,
    \sw_164_module_data_out[5] ,
    \sw_164_module_data_out[4] ,
    \sw_164_module_data_out[3] ,
    \sw_164_module_data_out[2] ,
    \sw_164_module_data_out[1] ,
    \sw_164_module_data_out[0] }));
 rc5_top rc5_top_043 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_043_module_data_in[7] ,
    \sw_043_module_data_in[6] ,
    \sw_043_module_data_in[5] ,
    \sw_043_module_data_in[4] ,
    \sw_043_module_data_in[3] ,
    \sw_043_module_data_in[2] ,
    \sw_043_module_data_in[1] ,
    \sw_043_module_data_in[0] }),
    .io_out({\sw_043_module_data_out[7] ,
    \sw_043_module_data_out[6] ,
    \sw_043_module_data_out[5] ,
    \sw_043_module_data_out[4] ,
    \sw_043_module_data_out[3] ,
    \sw_043_module_data_out[2] ,
    \sw_043_module_data_out[1] ,
    \sw_043_module_data_out[0] }));
 recepsaid_euclidean_algorithm recepsaid_euclidean_algorithm_133 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_133_module_data_in[7] ,
    \sw_133_module_data_in[6] ,
    \sw_133_module_data_in[5] ,
    \sw_133_module_data_in[4] ,
    \sw_133_module_data_in[3] ,
    \sw_133_module_data_in[2] ,
    \sw_133_module_data_in[1] ,
    \sw_133_module_data_in[0] }),
    .io_out({\sw_133_module_data_out[7] ,
    \sw_133_module_data_out[6] ,
    \sw_133_module_data_out[5] ,
    \sw_133_module_data_out[4] ,
    \sw_133_module_data_out[3] ,
    \sw_133_module_data_out[2] ,
    \sw_133_module_data_out[1] ,
    \sw_133_module_data_out[0] }));
 regymm_funnyblinky regymm_funnyblinky_098 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_098_module_data_in[7] ,
    \sw_098_module_data_in[6] ,
    \sw_098_module_data_in[5] ,
    \sw_098_module_data_in[4] ,
    \sw_098_module_data_in[3] ,
    \sw_098_module_data_in[2] ,
    \sw_098_module_data_in[1] ,
    \sw_098_module_data_in[0] }),
    .io_out({\sw_098_module_data_out[7] ,
    \sw_098_module_data_out[6] ,
    \sw_098_module_data_out[5] ,
    \sw_098_module_data_out[4] ,
    \sw_098_module_data_out[3] ,
    \sw_098_module_data_out[2] ,
    \sw_098_module_data_out[1] ,
    \sw_098_module_data_out[0] }));
 regymm_mcpi regymm_mcpi_097 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_097_module_data_in[7] ,
    \sw_097_module_data_in[6] ,
    \sw_097_module_data_in[5] ,
    \sw_097_module_data_in[4] ,
    \sw_097_module_data_in[3] ,
    \sw_097_module_data_in[2] ,
    \sw_097_module_data_in[1] ,
    \sw_097_module_data_in[0] }),
    .io_out({\sw_097_module_data_out[7] ,
    \sw_097_module_data_out[6] ,
    \sw_097_module_data_out[5] ,
    \sw_097_module_data_out[4] ,
    \sw_097_module_data_out[3] ,
    \sw_097_module_data_out[2] ,
    \sw_097_module_data_out[1] ,
    \sw_097_module_data_out[0] }));
 rglenn_hex_to_7_seg rglenn_hex_to_7_seg_121 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_121_module_data_in[7] ,
    \sw_121_module_data_in[6] ,
    \sw_121_module_data_in[5] ,
    \sw_121_module_data_in[4] ,
    \sw_121_module_data_in[3] ,
    \sw_121_module_data_in[2] ,
    \sw_121_module_data_in[1] ,
    \sw_121_module_data_in[0] }),
    .io_out({\sw_121_module_data_out[7] ,
    \sw_121_module_data_out[6] ,
    \sw_121_module_data_out[5] ,
    \sw_121_module_data_out[4] ,
    \sw_121_module_data_out[3] ,
    \sw_121_module_data_out[2] ,
    \sw_121_module_data_out[1] ,
    \sw_121_module_data_out[0] }));
 rolfmobile99_alu_fsm_top rolfmobile99_alu_fsm_top_035 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_035_module_data_in[7] ,
    \sw_035_module_data_in[6] ,
    \sw_035_module_data_in[5] ,
    \sw_035_module_data_in[4] ,
    \sw_035_module_data_in[3] ,
    \sw_035_module_data_in[2] ,
    \sw_035_module_data_in[1] ,
    \sw_035_module_data_in[0] }),
    .io_out({\sw_035_module_data_out[7] ,
    \sw_035_module_data_out[6] ,
    \sw_035_module_data_out[5] ,
    \sw_035_module_data_out[4] ,
    \sw_035_module_data_out[3] ,
    \sw_035_module_data_out[2] ,
    \sw_035_module_data_out[1] ,
    \sw_035_module_data_out[0] }));
 rotary_encoder rotary_encoder_113 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_113_module_data_in[7] ,
    \sw_113_module_data_in[6] ,
    \sw_113_module_data_in[5] ,
    \sw_113_module_data_in[4] ,
    \sw_113_module_data_in[3] ,
    \sw_113_module_data_in[2] ,
    \sw_113_module_data_in[1] ,
    \sw_113_module_data_in[0] }),
    .io_out({\sw_113_module_data_out[7] ,
    \sw_113_module_data_out[6] ,
    \sw_113_module_data_out[5] ,
    \sw_113_module_data_out[4] ,
    \sw_113_module_data_out[3] ,
    \sw_113_module_data_out[2] ,
    \sw_113_module_data_out[1] ,
    \sw_113_module_data_out[0] }));
 s4ga s4ga_006 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_006_module_data_in[7] ,
    \sw_006_module_data_in[6] ,
    \sw_006_module_data_in[5] ,
    \sw_006_module_data_in[4] ,
    \sw_006_module_data_in[3] ,
    \sw_006_module_data_in[2] ,
    \sw_006_module_data_in[1] ,
    \sw_006_module_data_in[0] }),
    .io_out({\sw_006_module_data_out[7] ,
    \sw_006_module_data_out[6] ,
    \sw_006_module_data_out[5] ,
    \sw_006_module_data_out[4] ,
    \sw_006_module_data_out[3] ,
    \sw_006_module_data_out[2] ,
    \sw_006_module_data_out[1] ,
    \sw_006_module_data_out[0] }));
 scan_controller scan_controller (.clk(wb_clk_i),
    .la_scan_clk_in(la_data_in[0]),
    .la_scan_data_in(la_data_in[1]),
    .la_scan_data_out(la_data_out[0]),
    .la_scan_latch_en(la_data_in[3]),
    .la_scan_select(la_data_in[2]),
    .ready(io_out[37]),
    .reset(wb_rst_i),
    .scan_clk_in(sc_clk_in),
    .scan_clk_out(sc_clk_out),
    .scan_data_in(sc_data_in),
    .scan_data_out(sc_data_out),
    .scan_latch_en(sc_latch_out),
    .scan_select(sc_scan_out),
    .set_clk_div(io_in[11]),
    .slow_clk(io_out[10]),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .active_select({io_in[20],
    io_in[19],
    io_in[18],
    io_in[17],
    io_in[16],
    io_in[15],
    io_in[14],
    io_in[13],
    io_in[12]}),
    .driver_sel({io_in[9],
    io_in[8]}),
    .inputs({io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21]}),
    .oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .outputs({io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29]}));
 scanchain scanchain_000 (.clk_in(sc_clk_out),
    .clk_out(sw_000_clk_out),
    .data_in(sc_data_out),
    .data_out(sw_000_data_out),
    .latch_enable_in(sc_latch_out),
    .latch_enable_out(sw_000_latch_out),
    .scan_select_in(sc_scan_out),
    .scan_select_out(sw_000_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_000_module_data_in[7] ,
    \sw_000_module_data_in[6] ,
    \sw_000_module_data_in[5] ,
    \sw_000_module_data_in[4] ,
    \sw_000_module_data_in[3] ,
    \sw_000_module_data_in[2] ,
    \sw_000_module_data_in[1] ,
    \sw_000_module_data_in[0] }),
    .module_data_out({\sw_000_module_data_out[7] ,
    \sw_000_module_data_out[6] ,
    \sw_000_module_data_out[5] ,
    \sw_000_module_data_out[4] ,
    \sw_000_module_data_out[3] ,
    \sw_000_module_data_out[2] ,
    \sw_000_module_data_out[1] ,
    \sw_000_module_data_out[0] }));
 scanchain scanchain_001 (.clk_in(sw_000_clk_out),
    .clk_out(sw_001_clk_out),
    .data_in(sw_000_data_out),
    .data_out(sw_001_data_out),
    .latch_enable_in(sw_000_latch_out),
    .latch_enable_out(sw_001_latch_out),
    .scan_select_in(sw_000_scan_out),
    .scan_select_out(sw_001_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_001_module_data_in[7] ,
    \sw_001_module_data_in[6] ,
    \sw_001_module_data_in[5] ,
    \sw_001_module_data_in[4] ,
    \sw_001_module_data_in[3] ,
    \sw_001_module_data_in[2] ,
    \sw_001_module_data_in[1] ,
    \sw_001_module_data_in[0] }),
    .module_data_out({\sw_001_module_data_out[7] ,
    \sw_001_module_data_out[6] ,
    \sw_001_module_data_out[5] ,
    \sw_001_module_data_out[4] ,
    \sw_001_module_data_out[3] ,
    \sw_001_module_data_out[2] ,
    \sw_001_module_data_out[1] ,
    \sw_001_module_data_out[0] }));
 scanchain scanchain_002 (.clk_in(sw_001_clk_out),
    .clk_out(sw_002_clk_out),
    .data_in(sw_001_data_out),
    .data_out(sw_002_data_out),
    .latch_enable_in(sw_001_latch_out),
    .latch_enable_out(sw_002_latch_out),
    .scan_select_in(sw_001_scan_out),
    .scan_select_out(sw_002_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_002_module_data_in[7] ,
    \sw_002_module_data_in[6] ,
    \sw_002_module_data_in[5] ,
    \sw_002_module_data_in[4] ,
    \sw_002_module_data_in[3] ,
    \sw_002_module_data_in[2] ,
    \sw_002_module_data_in[1] ,
    \sw_002_module_data_in[0] }),
    .module_data_out({\sw_002_module_data_out[7] ,
    \sw_002_module_data_out[6] ,
    \sw_002_module_data_out[5] ,
    \sw_002_module_data_out[4] ,
    \sw_002_module_data_out[3] ,
    \sw_002_module_data_out[2] ,
    \sw_002_module_data_out[1] ,
    \sw_002_module_data_out[0] }));
 scanchain scanchain_003 (.clk_in(sw_002_clk_out),
    .clk_out(sw_003_clk_out),
    .data_in(sw_002_data_out),
    .data_out(sw_003_data_out),
    .latch_enable_in(sw_002_latch_out),
    .latch_enable_out(sw_003_latch_out),
    .scan_select_in(sw_002_scan_out),
    .scan_select_out(sw_003_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_003_module_data_in[7] ,
    \sw_003_module_data_in[6] ,
    \sw_003_module_data_in[5] ,
    \sw_003_module_data_in[4] ,
    \sw_003_module_data_in[3] ,
    \sw_003_module_data_in[2] ,
    \sw_003_module_data_in[1] ,
    \sw_003_module_data_in[0] }),
    .module_data_out({\sw_003_module_data_out[7] ,
    \sw_003_module_data_out[6] ,
    \sw_003_module_data_out[5] ,
    \sw_003_module_data_out[4] ,
    \sw_003_module_data_out[3] ,
    \sw_003_module_data_out[2] ,
    \sw_003_module_data_out[1] ,
    \sw_003_module_data_out[0] }));
 scanchain scanchain_004 (.clk_in(sw_003_clk_out),
    .clk_out(sw_004_clk_out),
    .data_in(sw_003_data_out),
    .data_out(sw_004_data_out),
    .latch_enable_in(sw_003_latch_out),
    .latch_enable_out(sw_004_latch_out),
    .scan_select_in(sw_003_scan_out),
    .scan_select_out(sw_004_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_004_module_data_in[7] ,
    \sw_004_module_data_in[6] ,
    \sw_004_module_data_in[5] ,
    \sw_004_module_data_in[4] ,
    \sw_004_module_data_in[3] ,
    \sw_004_module_data_in[2] ,
    \sw_004_module_data_in[1] ,
    \sw_004_module_data_in[0] }),
    .module_data_out({\sw_004_module_data_out[7] ,
    \sw_004_module_data_out[6] ,
    \sw_004_module_data_out[5] ,
    \sw_004_module_data_out[4] ,
    \sw_004_module_data_out[3] ,
    \sw_004_module_data_out[2] ,
    \sw_004_module_data_out[1] ,
    \sw_004_module_data_out[0] }));
 scanchain scanchain_005 (.clk_in(sw_004_clk_out),
    .clk_out(sw_005_clk_out),
    .data_in(sw_004_data_out),
    .data_out(sw_005_data_out),
    .latch_enable_in(sw_004_latch_out),
    .latch_enable_out(sw_005_latch_out),
    .scan_select_in(sw_004_scan_out),
    .scan_select_out(sw_005_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_005_module_data_in[7] ,
    \sw_005_module_data_in[6] ,
    \sw_005_module_data_in[5] ,
    \sw_005_module_data_in[4] ,
    \sw_005_module_data_in[3] ,
    \sw_005_module_data_in[2] ,
    \sw_005_module_data_in[1] ,
    \sw_005_module_data_in[0] }),
    .module_data_out({\sw_005_module_data_out[7] ,
    \sw_005_module_data_out[6] ,
    \sw_005_module_data_out[5] ,
    \sw_005_module_data_out[4] ,
    \sw_005_module_data_out[3] ,
    \sw_005_module_data_out[2] ,
    \sw_005_module_data_out[1] ,
    \sw_005_module_data_out[0] }));
 scanchain scanchain_006 (.clk_in(sw_005_clk_out),
    .clk_out(sw_006_clk_out),
    .data_in(sw_005_data_out),
    .data_out(sw_006_data_out),
    .latch_enable_in(sw_005_latch_out),
    .latch_enable_out(sw_006_latch_out),
    .scan_select_in(sw_005_scan_out),
    .scan_select_out(sw_006_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_006_module_data_in[7] ,
    \sw_006_module_data_in[6] ,
    \sw_006_module_data_in[5] ,
    \sw_006_module_data_in[4] ,
    \sw_006_module_data_in[3] ,
    \sw_006_module_data_in[2] ,
    \sw_006_module_data_in[1] ,
    \sw_006_module_data_in[0] }),
    .module_data_out({\sw_006_module_data_out[7] ,
    \sw_006_module_data_out[6] ,
    \sw_006_module_data_out[5] ,
    \sw_006_module_data_out[4] ,
    \sw_006_module_data_out[3] ,
    \sw_006_module_data_out[2] ,
    \sw_006_module_data_out[1] ,
    \sw_006_module_data_out[0] }));
 scanchain scanchain_007 (.clk_in(sw_006_clk_out),
    .clk_out(sw_007_clk_out),
    .data_in(sw_006_data_out),
    .data_out(sw_007_data_out),
    .latch_enable_in(sw_006_latch_out),
    .latch_enable_out(sw_007_latch_out),
    .scan_select_in(sw_006_scan_out),
    .scan_select_out(sw_007_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_007_module_data_in[7] ,
    \sw_007_module_data_in[6] ,
    \sw_007_module_data_in[5] ,
    \sw_007_module_data_in[4] ,
    \sw_007_module_data_in[3] ,
    \sw_007_module_data_in[2] ,
    \sw_007_module_data_in[1] ,
    \sw_007_module_data_in[0] }),
    .module_data_out({\sw_007_module_data_out[7] ,
    \sw_007_module_data_out[6] ,
    \sw_007_module_data_out[5] ,
    \sw_007_module_data_out[4] ,
    \sw_007_module_data_out[3] ,
    \sw_007_module_data_out[2] ,
    \sw_007_module_data_out[1] ,
    \sw_007_module_data_out[0] }));
 scanchain scanchain_008 (.clk_in(sw_007_clk_out),
    .clk_out(sw_008_clk_out),
    .data_in(sw_007_data_out),
    .data_out(sw_008_data_out),
    .latch_enable_in(sw_007_latch_out),
    .latch_enable_out(sw_008_latch_out),
    .scan_select_in(sw_007_scan_out),
    .scan_select_out(sw_008_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_008_module_data_in[7] ,
    \sw_008_module_data_in[6] ,
    \sw_008_module_data_in[5] ,
    \sw_008_module_data_in[4] ,
    \sw_008_module_data_in[3] ,
    \sw_008_module_data_in[2] ,
    \sw_008_module_data_in[1] ,
    \sw_008_module_data_in[0] }),
    .module_data_out({\sw_008_module_data_out[7] ,
    \sw_008_module_data_out[6] ,
    \sw_008_module_data_out[5] ,
    \sw_008_module_data_out[4] ,
    \sw_008_module_data_out[3] ,
    \sw_008_module_data_out[2] ,
    \sw_008_module_data_out[1] ,
    \sw_008_module_data_out[0] }));
 scanchain scanchain_009 (.clk_in(sw_008_clk_out),
    .clk_out(sw_009_clk_out),
    .data_in(sw_008_data_out),
    .data_out(sw_009_data_out),
    .latch_enable_in(sw_008_latch_out),
    .latch_enable_out(sw_009_latch_out),
    .scan_select_in(sw_008_scan_out),
    .scan_select_out(sw_009_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_009_module_data_in[7] ,
    \sw_009_module_data_in[6] ,
    \sw_009_module_data_in[5] ,
    \sw_009_module_data_in[4] ,
    \sw_009_module_data_in[3] ,
    \sw_009_module_data_in[2] ,
    \sw_009_module_data_in[1] ,
    \sw_009_module_data_in[0] }),
    .module_data_out({\sw_009_module_data_out[7] ,
    \sw_009_module_data_out[6] ,
    \sw_009_module_data_out[5] ,
    \sw_009_module_data_out[4] ,
    \sw_009_module_data_out[3] ,
    \sw_009_module_data_out[2] ,
    \sw_009_module_data_out[1] ,
    \sw_009_module_data_out[0] }));
 scanchain scanchain_010 (.clk_in(sw_009_clk_out),
    .clk_out(sw_010_clk_out),
    .data_in(sw_009_data_out),
    .data_out(sw_010_data_out),
    .latch_enable_in(sw_009_latch_out),
    .latch_enable_out(sw_010_latch_out),
    .scan_select_in(sw_009_scan_out),
    .scan_select_out(sw_010_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_010_module_data_in[7] ,
    \sw_010_module_data_in[6] ,
    \sw_010_module_data_in[5] ,
    \sw_010_module_data_in[4] ,
    \sw_010_module_data_in[3] ,
    \sw_010_module_data_in[2] ,
    \sw_010_module_data_in[1] ,
    \sw_010_module_data_in[0] }),
    .module_data_out({\sw_010_module_data_out[7] ,
    \sw_010_module_data_out[6] ,
    \sw_010_module_data_out[5] ,
    \sw_010_module_data_out[4] ,
    \sw_010_module_data_out[3] ,
    \sw_010_module_data_out[2] ,
    \sw_010_module_data_out[1] ,
    \sw_010_module_data_out[0] }));
 scanchain scanchain_011 (.clk_in(sw_010_clk_out),
    .clk_out(sw_011_clk_out),
    .data_in(sw_010_data_out),
    .data_out(sw_011_data_out),
    .latch_enable_in(sw_010_latch_out),
    .latch_enable_out(sw_011_latch_out),
    .scan_select_in(sw_010_scan_out),
    .scan_select_out(sw_011_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_011_module_data_in[7] ,
    \sw_011_module_data_in[6] ,
    \sw_011_module_data_in[5] ,
    \sw_011_module_data_in[4] ,
    \sw_011_module_data_in[3] ,
    \sw_011_module_data_in[2] ,
    \sw_011_module_data_in[1] ,
    \sw_011_module_data_in[0] }),
    .module_data_out({\sw_011_module_data_out[7] ,
    \sw_011_module_data_out[6] ,
    \sw_011_module_data_out[5] ,
    \sw_011_module_data_out[4] ,
    \sw_011_module_data_out[3] ,
    \sw_011_module_data_out[2] ,
    \sw_011_module_data_out[1] ,
    \sw_011_module_data_out[0] }));
 scanchain scanchain_012 (.clk_in(sw_011_clk_out),
    .clk_out(sw_012_clk_out),
    .data_in(sw_011_data_out),
    .data_out(sw_012_data_out),
    .latch_enable_in(sw_011_latch_out),
    .latch_enable_out(sw_012_latch_out),
    .scan_select_in(sw_011_scan_out),
    .scan_select_out(sw_012_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_012_module_data_in[7] ,
    \sw_012_module_data_in[6] ,
    \sw_012_module_data_in[5] ,
    \sw_012_module_data_in[4] ,
    \sw_012_module_data_in[3] ,
    \sw_012_module_data_in[2] ,
    \sw_012_module_data_in[1] ,
    \sw_012_module_data_in[0] }),
    .module_data_out({\sw_012_module_data_out[7] ,
    \sw_012_module_data_out[6] ,
    \sw_012_module_data_out[5] ,
    \sw_012_module_data_out[4] ,
    \sw_012_module_data_out[3] ,
    \sw_012_module_data_out[2] ,
    \sw_012_module_data_out[1] ,
    \sw_012_module_data_out[0] }));
 scanchain scanchain_013 (.clk_in(sw_012_clk_out),
    .clk_out(sw_013_clk_out),
    .data_in(sw_012_data_out),
    .data_out(sw_013_data_out),
    .latch_enable_in(sw_012_latch_out),
    .latch_enable_out(sw_013_latch_out),
    .scan_select_in(sw_012_scan_out),
    .scan_select_out(sw_013_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_013_module_data_in[7] ,
    \sw_013_module_data_in[6] ,
    \sw_013_module_data_in[5] ,
    \sw_013_module_data_in[4] ,
    \sw_013_module_data_in[3] ,
    \sw_013_module_data_in[2] ,
    \sw_013_module_data_in[1] ,
    \sw_013_module_data_in[0] }),
    .module_data_out({\sw_013_module_data_out[7] ,
    \sw_013_module_data_out[6] ,
    \sw_013_module_data_out[5] ,
    \sw_013_module_data_out[4] ,
    \sw_013_module_data_out[3] ,
    \sw_013_module_data_out[2] ,
    \sw_013_module_data_out[1] ,
    \sw_013_module_data_out[0] }));
 scanchain scanchain_014 (.clk_in(sw_013_clk_out),
    .clk_out(sw_014_clk_out),
    .data_in(sw_013_data_out),
    .data_out(sw_014_data_out),
    .latch_enable_in(sw_013_latch_out),
    .latch_enable_out(sw_014_latch_out),
    .scan_select_in(sw_013_scan_out),
    .scan_select_out(sw_014_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_014_module_data_in[7] ,
    \sw_014_module_data_in[6] ,
    \sw_014_module_data_in[5] ,
    \sw_014_module_data_in[4] ,
    \sw_014_module_data_in[3] ,
    \sw_014_module_data_in[2] ,
    \sw_014_module_data_in[1] ,
    \sw_014_module_data_in[0] }),
    .module_data_out({\sw_014_module_data_out[7] ,
    \sw_014_module_data_out[6] ,
    \sw_014_module_data_out[5] ,
    \sw_014_module_data_out[4] ,
    \sw_014_module_data_out[3] ,
    \sw_014_module_data_out[2] ,
    \sw_014_module_data_out[1] ,
    \sw_014_module_data_out[0] }));
 scanchain scanchain_015 (.clk_in(sw_014_clk_out),
    .clk_out(sw_015_clk_out),
    .data_in(sw_014_data_out),
    .data_out(sw_015_data_out),
    .latch_enable_in(sw_014_latch_out),
    .latch_enable_out(sw_015_latch_out),
    .scan_select_in(sw_014_scan_out),
    .scan_select_out(sw_015_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_015_module_data_in[7] ,
    \sw_015_module_data_in[6] ,
    \sw_015_module_data_in[5] ,
    \sw_015_module_data_in[4] ,
    \sw_015_module_data_in[3] ,
    \sw_015_module_data_in[2] ,
    \sw_015_module_data_in[1] ,
    \sw_015_module_data_in[0] }),
    .module_data_out({\sw_015_module_data_out[7] ,
    \sw_015_module_data_out[6] ,
    \sw_015_module_data_out[5] ,
    \sw_015_module_data_out[4] ,
    \sw_015_module_data_out[3] ,
    \sw_015_module_data_out[2] ,
    \sw_015_module_data_out[1] ,
    \sw_015_module_data_out[0] }));
 scanchain scanchain_016 (.clk_in(sw_015_clk_out),
    .clk_out(sw_016_clk_out),
    .data_in(sw_015_data_out),
    .data_out(sw_016_data_out),
    .latch_enable_in(sw_015_latch_out),
    .latch_enable_out(sw_016_latch_out),
    .scan_select_in(sw_015_scan_out),
    .scan_select_out(sw_016_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_016_module_data_in[7] ,
    \sw_016_module_data_in[6] ,
    \sw_016_module_data_in[5] ,
    \sw_016_module_data_in[4] ,
    \sw_016_module_data_in[3] ,
    \sw_016_module_data_in[2] ,
    \sw_016_module_data_in[1] ,
    \sw_016_module_data_in[0] }),
    .module_data_out({\sw_016_module_data_out[7] ,
    \sw_016_module_data_out[6] ,
    \sw_016_module_data_out[5] ,
    \sw_016_module_data_out[4] ,
    \sw_016_module_data_out[3] ,
    \sw_016_module_data_out[2] ,
    \sw_016_module_data_out[1] ,
    \sw_016_module_data_out[0] }));
 scanchain scanchain_017 (.clk_in(sw_016_clk_out),
    .clk_out(sw_017_clk_out),
    .data_in(sw_016_data_out),
    .data_out(sw_017_data_out),
    .latch_enable_in(sw_016_latch_out),
    .latch_enable_out(sw_017_latch_out),
    .scan_select_in(sw_016_scan_out),
    .scan_select_out(sw_017_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_017_module_data_in[7] ,
    \sw_017_module_data_in[6] ,
    \sw_017_module_data_in[5] ,
    \sw_017_module_data_in[4] ,
    \sw_017_module_data_in[3] ,
    \sw_017_module_data_in[2] ,
    \sw_017_module_data_in[1] ,
    \sw_017_module_data_in[0] }),
    .module_data_out({\sw_017_module_data_out[7] ,
    \sw_017_module_data_out[6] ,
    \sw_017_module_data_out[5] ,
    \sw_017_module_data_out[4] ,
    \sw_017_module_data_out[3] ,
    \sw_017_module_data_out[2] ,
    \sw_017_module_data_out[1] ,
    \sw_017_module_data_out[0] }));
 scanchain scanchain_018 (.clk_in(sw_017_clk_out),
    .clk_out(sw_018_clk_out),
    .data_in(sw_017_data_out),
    .data_out(sw_018_data_out),
    .latch_enable_in(sw_017_latch_out),
    .latch_enable_out(sw_018_latch_out),
    .scan_select_in(sw_017_scan_out),
    .scan_select_out(sw_018_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_018_module_data_in[7] ,
    \sw_018_module_data_in[6] ,
    \sw_018_module_data_in[5] ,
    \sw_018_module_data_in[4] ,
    \sw_018_module_data_in[3] ,
    \sw_018_module_data_in[2] ,
    \sw_018_module_data_in[1] ,
    \sw_018_module_data_in[0] }),
    .module_data_out({\sw_018_module_data_out[7] ,
    \sw_018_module_data_out[6] ,
    \sw_018_module_data_out[5] ,
    \sw_018_module_data_out[4] ,
    \sw_018_module_data_out[3] ,
    \sw_018_module_data_out[2] ,
    \sw_018_module_data_out[1] ,
    \sw_018_module_data_out[0] }));
 scanchain scanchain_019 (.clk_in(sw_018_clk_out),
    .clk_out(sw_019_clk_out),
    .data_in(sw_018_data_out),
    .data_out(sw_019_data_out),
    .latch_enable_in(sw_018_latch_out),
    .latch_enable_out(sw_019_latch_out),
    .scan_select_in(sw_018_scan_out),
    .scan_select_out(sw_019_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_019_module_data_in[7] ,
    \sw_019_module_data_in[6] ,
    \sw_019_module_data_in[5] ,
    \sw_019_module_data_in[4] ,
    \sw_019_module_data_in[3] ,
    \sw_019_module_data_in[2] ,
    \sw_019_module_data_in[1] ,
    \sw_019_module_data_in[0] }),
    .module_data_out({\sw_019_module_data_out[7] ,
    \sw_019_module_data_out[6] ,
    \sw_019_module_data_out[5] ,
    \sw_019_module_data_out[4] ,
    \sw_019_module_data_out[3] ,
    \sw_019_module_data_out[2] ,
    \sw_019_module_data_out[1] ,
    \sw_019_module_data_out[0] }));
 scanchain scanchain_020 (.clk_in(sw_019_clk_out),
    .clk_out(sw_020_clk_out),
    .data_in(sw_019_data_out),
    .data_out(sw_020_data_out),
    .latch_enable_in(sw_019_latch_out),
    .latch_enable_out(sw_020_latch_out),
    .scan_select_in(sw_019_scan_out),
    .scan_select_out(sw_020_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_020_module_data_in[7] ,
    \sw_020_module_data_in[6] ,
    \sw_020_module_data_in[5] ,
    \sw_020_module_data_in[4] ,
    \sw_020_module_data_in[3] ,
    \sw_020_module_data_in[2] ,
    \sw_020_module_data_in[1] ,
    \sw_020_module_data_in[0] }),
    .module_data_out({\sw_020_module_data_out[7] ,
    \sw_020_module_data_out[6] ,
    \sw_020_module_data_out[5] ,
    \sw_020_module_data_out[4] ,
    \sw_020_module_data_out[3] ,
    \sw_020_module_data_out[2] ,
    \sw_020_module_data_out[1] ,
    \sw_020_module_data_out[0] }));
 scanchain scanchain_021 (.clk_in(sw_020_clk_out),
    .clk_out(sw_021_clk_out),
    .data_in(sw_020_data_out),
    .data_out(sw_021_data_out),
    .latch_enable_in(sw_020_latch_out),
    .latch_enable_out(sw_021_latch_out),
    .scan_select_in(sw_020_scan_out),
    .scan_select_out(sw_021_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_021_module_data_in[7] ,
    \sw_021_module_data_in[6] ,
    \sw_021_module_data_in[5] ,
    \sw_021_module_data_in[4] ,
    \sw_021_module_data_in[3] ,
    \sw_021_module_data_in[2] ,
    \sw_021_module_data_in[1] ,
    \sw_021_module_data_in[0] }),
    .module_data_out({\sw_021_module_data_out[7] ,
    \sw_021_module_data_out[6] ,
    \sw_021_module_data_out[5] ,
    \sw_021_module_data_out[4] ,
    \sw_021_module_data_out[3] ,
    \sw_021_module_data_out[2] ,
    \sw_021_module_data_out[1] ,
    \sw_021_module_data_out[0] }));
 scanchain scanchain_022 (.clk_in(sw_021_clk_out),
    .clk_out(sw_022_clk_out),
    .data_in(sw_021_data_out),
    .data_out(sw_022_data_out),
    .latch_enable_in(sw_021_latch_out),
    .latch_enable_out(sw_022_latch_out),
    .scan_select_in(sw_021_scan_out),
    .scan_select_out(sw_022_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_022_module_data_in[7] ,
    \sw_022_module_data_in[6] ,
    \sw_022_module_data_in[5] ,
    \sw_022_module_data_in[4] ,
    \sw_022_module_data_in[3] ,
    \sw_022_module_data_in[2] ,
    \sw_022_module_data_in[1] ,
    \sw_022_module_data_in[0] }),
    .module_data_out({\sw_022_module_data_out[7] ,
    \sw_022_module_data_out[6] ,
    \sw_022_module_data_out[5] ,
    \sw_022_module_data_out[4] ,
    \sw_022_module_data_out[3] ,
    \sw_022_module_data_out[2] ,
    \sw_022_module_data_out[1] ,
    \sw_022_module_data_out[0] }));
 scanchain scanchain_023 (.clk_in(sw_022_clk_out),
    .clk_out(sw_023_clk_out),
    .data_in(sw_022_data_out),
    .data_out(sw_023_data_out),
    .latch_enable_in(sw_022_latch_out),
    .latch_enable_out(sw_023_latch_out),
    .scan_select_in(sw_022_scan_out),
    .scan_select_out(sw_023_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_023_module_data_in[7] ,
    \sw_023_module_data_in[6] ,
    \sw_023_module_data_in[5] ,
    \sw_023_module_data_in[4] ,
    \sw_023_module_data_in[3] ,
    \sw_023_module_data_in[2] ,
    \sw_023_module_data_in[1] ,
    \sw_023_module_data_in[0] }),
    .module_data_out({\sw_023_module_data_out[7] ,
    \sw_023_module_data_out[6] ,
    \sw_023_module_data_out[5] ,
    \sw_023_module_data_out[4] ,
    \sw_023_module_data_out[3] ,
    \sw_023_module_data_out[2] ,
    \sw_023_module_data_out[1] ,
    \sw_023_module_data_out[0] }));
 scanchain scanchain_024 (.clk_in(sw_023_clk_out),
    .clk_out(sw_024_clk_out),
    .data_in(sw_023_data_out),
    .data_out(sw_024_data_out),
    .latch_enable_in(sw_023_latch_out),
    .latch_enable_out(sw_024_latch_out),
    .scan_select_in(sw_023_scan_out),
    .scan_select_out(sw_024_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_024_module_data_in[7] ,
    \sw_024_module_data_in[6] ,
    \sw_024_module_data_in[5] ,
    \sw_024_module_data_in[4] ,
    \sw_024_module_data_in[3] ,
    \sw_024_module_data_in[2] ,
    \sw_024_module_data_in[1] ,
    \sw_024_module_data_in[0] }),
    .module_data_out({\sw_024_module_data_out[7] ,
    \sw_024_module_data_out[6] ,
    \sw_024_module_data_out[5] ,
    \sw_024_module_data_out[4] ,
    \sw_024_module_data_out[3] ,
    \sw_024_module_data_out[2] ,
    \sw_024_module_data_out[1] ,
    \sw_024_module_data_out[0] }));
 scanchain scanchain_025 (.clk_in(sw_024_clk_out),
    .clk_out(sw_025_clk_out),
    .data_in(sw_024_data_out),
    .data_out(sw_025_data_out),
    .latch_enable_in(sw_024_latch_out),
    .latch_enable_out(sw_025_latch_out),
    .scan_select_in(sw_024_scan_out),
    .scan_select_out(sw_025_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_025_module_data_in[7] ,
    \sw_025_module_data_in[6] ,
    \sw_025_module_data_in[5] ,
    \sw_025_module_data_in[4] ,
    \sw_025_module_data_in[3] ,
    \sw_025_module_data_in[2] ,
    \sw_025_module_data_in[1] ,
    \sw_025_module_data_in[0] }),
    .module_data_out({\sw_025_module_data_out[7] ,
    \sw_025_module_data_out[6] ,
    \sw_025_module_data_out[5] ,
    \sw_025_module_data_out[4] ,
    \sw_025_module_data_out[3] ,
    \sw_025_module_data_out[2] ,
    \sw_025_module_data_out[1] ,
    \sw_025_module_data_out[0] }));
 scanchain scanchain_026 (.clk_in(sw_025_clk_out),
    .clk_out(sw_026_clk_out),
    .data_in(sw_025_data_out),
    .data_out(sw_026_data_out),
    .latch_enable_in(sw_025_latch_out),
    .latch_enable_out(sw_026_latch_out),
    .scan_select_in(sw_025_scan_out),
    .scan_select_out(sw_026_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_026_module_data_in[7] ,
    \sw_026_module_data_in[6] ,
    \sw_026_module_data_in[5] ,
    \sw_026_module_data_in[4] ,
    \sw_026_module_data_in[3] ,
    \sw_026_module_data_in[2] ,
    \sw_026_module_data_in[1] ,
    \sw_026_module_data_in[0] }),
    .module_data_out({\sw_026_module_data_out[7] ,
    \sw_026_module_data_out[6] ,
    \sw_026_module_data_out[5] ,
    \sw_026_module_data_out[4] ,
    \sw_026_module_data_out[3] ,
    \sw_026_module_data_out[2] ,
    \sw_026_module_data_out[1] ,
    \sw_026_module_data_out[0] }));
 scanchain scanchain_027 (.clk_in(sw_026_clk_out),
    .clk_out(sw_027_clk_out),
    .data_in(sw_026_data_out),
    .data_out(sw_027_data_out),
    .latch_enable_in(sw_026_latch_out),
    .latch_enable_out(sw_027_latch_out),
    .scan_select_in(sw_026_scan_out),
    .scan_select_out(sw_027_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_027_module_data_in[7] ,
    \sw_027_module_data_in[6] ,
    \sw_027_module_data_in[5] ,
    \sw_027_module_data_in[4] ,
    \sw_027_module_data_in[3] ,
    \sw_027_module_data_in[2] ,
    \sw_027_module_data_in[1] ,
    \sw_027_module_data_in[0] }),
    .module_data_out({\sw_027_module_data_out[7] ,
    \sw_027_module_data_out[6] ,
    \sw_027_module_data_out[5] ,
    \sw_027_module_data_out[4] ,
    \sw_027_module_data_out[3] ,
    \sw_027_module_data_out[2] ,
    \sw_027_module_data_out[1] ,
    \sw_027_module_data_out[0] }));
 scanchain scanchain_028 (.clk_in(sw_027_clk_out),
    .clk_out(sw_028_clk_out),
    .data_in(sw_027_data_out),
    .data_out(sw_028_data_out),
    .latch_enable_in(sw_027_latch_out),
    .latch_enable_out(sw_028_latch_out),
    .scan_select_in(sw_027_scan_out),
    .scan_select_out(sw_028_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_028_module_data_in[7] ,
    \sw_028_module_data_in[6] ,
    \sw_028_module_data_in[5] ,
    \sw_028_module_data_in[4] ,
    \sw_028_module_data_in[3] ,
    \sw_028_module_data_in[2] ,
    \sw_028_module_data_in[1] ,
    \sw_028_module_data_in[0] }),
    .module_data_out({\sw_028_module_data_out[7] ,
    \sw_028_module_data_out[6] ,
    \sw_028_module_data_out[5] ,
    \sw_028_module_data_out[4] ,
    \sw_028_module_data_out[3] ,
    \sw_028_module_data_out[2] ,
    \sw_028_module_data_out[1] ,
    \sw_028_module_data_out[0] }));
 scanchain scanchain_029 (.clk_in(sw_028_clk_out),
    .clk_out(sw_029_clk_out),
    .data_in(sw_028_data_out),
    .data_out(sw_029_data_out),
    .latch_enable_in(sw_028_latch_out),
    .latch_enable_out(sw_029_latch_out),
    .scan_select_in(sw_028_scan_out),
    .scan_select_out(sw_029_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_029_module_data_in[7] ,
    \sw_029_module_data_in[6] ,
    \sw_029_module_data_in[5] ,
    \sw_029_module_data_in[4] ,
    \sw_029_module_data_in[3] ,
    \sw_029_module_data_in[2] ,
    \sw_029_module_data_in[1] ,
    \sw_029_module_data_in[0] }),
    .module_data_out({\sw_029_module_data_out[7] ,
    \sw_029_module_data_out[6] ,
    \sw_029_module_data_out[5] ,
    \sw_029_module_data_out[4] ,
    \sw_029_module_data_out[3] ,
    \sw_029_module_data_out[2] ,
    \sw_029_module_data_out[1] ,
    \sw_029_module_data_out[0] }));
 scanchain scanchain_030 (.clk_in(sw_029_clk_out),
    .clk_out(sw_030_clk_out),
    .data_in(sw_029_data_out),
    .data_out(sw_030_data_out),
    .latch_enable_in(sw_029_latch_out),
    .latch_enable_out(sw_030_latch_out),
    .scan_select_in(sw_029_scan_out),
    .scan_select_out(sw_030_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_030_module_data_in[7] ,
    \sw_030_module_data_in[6] ,
    \sw_030_module_data_in[5] ,
    \sw_030_module_data_in[4] ,
    \sw_030_module_data_in[3] ,
    \sw_030_module_data_in[2] ,
    \sw_030_module_data_in[1] ,
    \sw_030_module_data_in[0] }),
    .module_data_out({\sw_030_module_data_out[7] ,
    \sw_030_module_data_out[6] ,
    \sw_030_module_data_out[5] ,
    \sw_030_module_data_out[4] ,
    \sw_030_module_data_out[3] ,
    \sw_030_module_data_out[2] ,
    \sw_030_module_data_out[1] ,
    \sw_030_module_data_out[0] }));
 scanchain scanchain_031 (.clk_in(sw_030_clk_out),
    .clk_out(sw_031_clk_out),
    .data_in(sw_030_data_out),
    .data_out(sw_031_data_out),
    .latch_enable_in(sw_030_latch_out),
    .latch_enable_out(sw_031_latch_out),
    .scan_select_in(sw_030_scan_out),
    .scan_select_out(sw_031_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_031_module_data_in[7] ,
    \sw_031_module_data_in[6] ,
    \sw_031_module_data_in[5] ,
    \sw_031_module_data_in[4] ,
    \sw_031_module_data_in[3] ,
    \sw_031_module_data_in[2] ,
    \sw_031_module_data_in[1] ,
    \sw_031_module_data_in[0] }),
    .module_data_out({\sw_031_module_data_out[7] ,
    \sw_031_module_data_out[6] ,
    \sw_031_module_data_out[5] ,
    \sw_031_module_data_out[4] ,
    \sw_031_module_data_out[3] ,
    \sw_031_module_data_out[2] ,
    \sw_031_module_data_out[1] ,
    \sw_031_module_data_out[0] }));
 scanchain scanchain_032 (.clk_in(sw_031_clk_out),
    .clk_out(sw_032_clk_out),
    .data_in(sw_031_data_out),
    .data_out(sw_032_data_out),
    .latch_enable_in(sw_031_latch_out),
    .latch_enable_out(sw_032_latch_out),
    .scan_select_in(sw_031_scan_out),
    .scan_select_out(sw_032_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_032_module_data_in[7] ,
    \sw_032_module_data_in[6] ,
    \sw_032_module_data_in[5] ,
    \sw_032_module_data_in[4] ,
    \sw_032_module_data_in[3] ,
    \sw_032_module_data_in[2] ,
    \sw_032_module_data_in[1] ,
    \sw_032_module_data_in[0] }),
    .module_data_out({\sw_032_module_data_out[7] ,
    \sw_032_module_data_out[6] ,
    \sw_032_module_data_out[5] ,
    \sw_032_module_data_out[4] ,
    \sw_032_module_data_out[3] ,
    \sw_032_module_data_out[2] ,
    \sw_032_module_data_out[1] ,
    \sw_032_module_data_out[0] }));
 scanchain scanchain_033 (.clk_in(sw_032_clk_out),
    .clk_out(sw_033_clk_out),
    .data_in(sw_032_data_out),
    .data_out(sw_033_data_out),
    .latch_enable_in(sw_032_latch_out),
    .latch_enable_out(sw_033_latch_out),
    .scan_select_in(sw_032_scan_out),
    .scan_select_out(sw_033_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_033_module_data_in[7] ,
    \sw_033_module_data_in[6] ,
    \sw_033_module_data_in[5] ,
    \sw_033_module_data_in[4] ,
    \sw_033_module_data_in[3] ,
    \sw_033_module_data_in[2] ,
    \sw_033_module_data_in[1] ,
    \sw_033_module_data_in[0] }),
    .module_data_out({\sw_033_module_data_out[7] ,
    \sw_033_module_data_out[6] ,
    \sw_033_module_data_out[5] ,
    \sw_033_module_data_out[4] ,
    \sw_033_module_data_out[3] ,
    \sw_033_module_data_out[2] ,
    \sw_033_module_data_out[1] ,
    \sw_033_module_data_out[0] }));
 scanchain scanchain_034 (.clk_in(sw_033_clk_out),
    .clk_out(sw_034_clk_out),
    .data_in(sw_033_data_out),
    .data_out(sw_034_data_out),
    .latch_enable_in(sw_033_latch_out),
    .latch_enable_out(sw_034_latch_out),
    .scan_select_in(sw_033_scan_out),
    .scan_select_out(sw_034_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_034_module_data_in[7] ,
    \sw_034_module_data_in[6] ,
    \sw_034_module_data_in[5] ,
    \sw_034_module_data_in[4] ,
    \sw_034_module_data_in[3] ,
    \sw_034_module_data_in[2] ,
    \sw_034_module_data_in[1] ,
    \sw_034_module_data_in[0] }),
    .module_data_out({\sw_034_module_data_out[7] ,
    \sw_034_module_data_out[6] ,
    \sw_034_module_data_out[5] ,
    \sw_034_module_data_out[4] ,
    \sw_034_module_data_out[3] ,
    \sw_034_module_data_out[2] ,
    \sw_034_module_data_out[1] ,
    \sw_034_module_data_out[0] }));
 scanchain scanchain_035 (.clk_in(sw_034_clk_out),
    .clk_out(sw_035_clk_out),
    .data_in(sw_034_data_out),
    .data_out(sw_035_data_out),
    .latch_enable_in(sw_034_latch_out),
    .latch_enable_out(sw_035_latch_out),
    .scan_select_in(sw_034_scan_out),
    .scan_select_out(sw_035_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_035_module_data_in[7] ,
    \sw_035_module_data_in[6] ,
    \sw_035_module_data_in[5] ,
    \sw_035_module_data_in[4] ,
    \sw_035_module_data_in[3] ,
    \sw_035_module_data_in[2] ,
    \sw_035_module_data_in[1] ,
    \sw_035_module_data_in[0] }),
    .module_data_out({\sw_035_module_data_out[7] ,
    \sw_035_module_data_out[6] ,
    \sw_035_module_data_out[5] ,
    \sw_035_module_data_out[4] ,
    \sw_035_module_data_out[3] ,
    \sw_035_module_data_out[2] ,
    \sw_035_module_data_out[1] ,
    \sw_035_module_data_out[0] }));
 scanchain scanchain_036 (.clk_in(sw_035_clk_out),
    .clk_out(sw_036_clk_out),
    .data_in(sw_035_data_out),
    .data_out(sw_036_data_out),
    .latch_enable_in(sw_035_latch_out),
    .latch_enable_out(sw_036_latch_out),
    .scan_select_in(sw_035_scan_out),
    .scan_select_out(sw_036_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_036_module_data_in[7] ,
    \sw_036_module_data_in[6] ,
    \sw_036_module_data_in[5] ,
    \sw_036_module_data_in[4] ,
    \sw_036_module_data_in[3] ,
    \sw_036_module_data_in[2] ,
    \sw_036_module_data_in[1] ,
    \sw_036_module_data_in[0] }),
    .module_data_out({\sw_036_module_data_out[7] ,
    \sw_036_module_data_out[6] ,
    \sw_036_module_data_out[5] ,
    \sw_036_module_data_out[4] ,
    \sw_036_module_data_out[3] ,
    \sw_036_module_data_out[2] ,
    \sw_036_module_data_out[1] ,
    \sw_036_module_data_out[0] }));
 scanchain scanchain_037 (.clk_in(sw_036_clk_out),
    .clk_out(sw_037_clk_out),
    .data_in(sw_036_data_out),
    .data_out(sw_037_data_out),
    .latch_enable_in(sw_036_latch_out),
    .latch_enable_out(sw_037_latch_out),
    .scan_select_in(sw_036_scan_out),
    .scan_select_out(sw_037_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_037_module_data_in[7] ,
    \sw_037_module_data_in[6] ,
    \sw_037_module_data_in[5] ,
    \sw_037_module_data_in[4] ,
    \sw_037_module_data_in[3] ,
    \sw_037_module_data_in[2] ,
    \sw_037_module_data_in[1] ,
    \sw_037_module_data_in[0] }),
    .module_data_out({\sw_037_module_data_out[7] ,
    \sw_037_module_data_out[6] ,
    \sw_037_module_data_out[5] ,
    \sw_037_module_data_out[4] ,
    \sw_037_module_data_out[3] ,
    \sw_037_module_data_out[2] ,
    \sw_037_module_data_out[1] ,
    \sw_037_module_data_out[0] }));
 scanchain scanchain_038 (.clk_in(sw_037_clk_out),
    .clk_out(sw_038_clk_out),
    .data_in(sw_037_data_out),
    .data_out(sw_038_data_out),
    .latch_enable_in(sw_037_latch_out),
    .latch_enable_out(sw_038_latch_out),
    .scan_select_in(sw_037_scan_out),
    .scan_select_out(sw_038_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_038_module_data_in[7] ,
    \sw_038_module_data_in[6] ,
    \sw_038_module_data_in[5] ,
    \sw_038_module_data_in[4] ,
    \sw_038_module_data_in[3] ,
    \sw_038_module_data_in[2] ,
    \sw_038_module_data_in[1] ,
    \sw_038_module_data_in[0] }),
    .module_data_out({\sw_038_module_data_out[7] ,
    \sw_038_module_data_out[6] ,
    \sw_038_module_data_out[5] ,
    \sw_038_module_data_out[4] ,
    \sw_038_module_data_out[3] ,
    \sw_038_module_data_out[2] ,
    \sw_038_module_data_out[1] ,
    \sw_038_module_data_out[0] }));
 scanchain scanchain_039 (.clk_in(sw_038_clk_out),
    .clk_out(sw_039_clk_out),
    .data_in(sw_038_data_out),
    .data_out(sw_039_data_out),
    .latch_enable_in(sw_038_latch_out),
    .latch_enable_out(sw_039_latch_out),
    .scan_select_in(sw_038_scan_out),
    .scan_select_out(sw_039_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_039_module_data_in[7] ,
    \sw_039_module_data_in[6] ,
    \sw_039_module_data_in[5] ,
    \sw_039_module_data_in[4] ,
    \sw_039_module_data_in[3] ,
    \sw_039_module_data_in[2] ,
    \sw_039_module_data_in[1] ,
    \sw_039_module_data_in[0] }),
    .module_data_out({\sw_039_module_data_out[7] ,
    \sw_039_module_data_out[6] ,
    \sw_039_module_data_out[5] ,
    \sw_039_module_data_out[4] ,
    \sw_039_module_data_out[3] ,
    \sw_039_module_data_out[2] ,
    \sw_039_module_data_out[1] ,
    \sw_039_module_data_out[0] }));
 scanchain scanchain_040 (.clk_in(sw_039_clk_out),
    .clk_out(sw_040_clk_out),
    .data_in(sw_039_data_out),
    .data_out(sw_040_data_out),
    .latch_enable_in(sw_039_latch_out),
    .latch_enable_out(sw_040_latch_out),
    .scan_select_in(sw_039_scan_out),
    .scan_select_out(sw_040_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_040_module_data_in[7] ,
    \sw_040_module_data_in[6] ,
    \sw_040_module_data_in[5] ,
    \sw_040_module_data_in[4] ,
    \sw_040_module_data_in[3] ,
    \sw_040_module_data_in[2] ,
    \sw_040_module_data_in[1] ,
    \sw_040_module_data_in[0] }),
    .module_data_out({\sw_040_module_data_out[7] ,
    \sw_040_module_data_out[6] ,
    \sw_040_module_data_out[5] ,
    \sw_040_module_data_out[4] ,
    \sw_040_module_data_out[3] ,
    \sw_040_module_data_out[2] ,
    \sw_040_module_data_out[1] ,
    \sw_040_module_data_out[0] }));
 scanchain scanchain_041 (.clk_in(sw_040_clk_out),
    .clk_out(sw_041_clk_out),
    .data_in(sw_040_data_out),
    .data_out(sw_041_data_out),
    .latch_enable_in(sw_040_latch_out),
    .latch_enable_out(sw_041_latch_out),
    .scan_select_in(sw_040_scan_out),
    .scan_select_out(sw_041_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_041_module_data_in[7] ,
    \sw_041_module_data_in[6] ,
    \sw_041_module_data_in[5] ,
    \sw_041_module_data_in[4] ,
    \sw_041_module_data_in[3] ,
    \sw_041_module_data_in[2] ,
    \sw_041_module_data_in[1] ,
    \sw_041_module_data_in[0] }),
    .module_data_out({\sw_041_module_data_out[7] ,
    \sw_041_module_data_out[6] ,
    \sw_041_module_data_out[5] ,
    \sw_041_module_data_out[4] ,
    \sw_041_module_data_out[3] ,
    \sw_041_module_data_out[2] ,
    \sw_041_module_data_out[1] ,
    \sw_041_module_data_out[0] }));
 scanchain scanchain_042 (.clk_in(sw_041_clk_out),
    .clk_out(sw_042_clk_out),
    .data_in(sw_041_data_out),
    .data_out(sw_042_data_out),
    .latch_enable_in(sw_041_latch_out),
    .latch_enable_out(sw_042_latch_out),
    .scan_select_in(sw_041_scan_out),
    .scan_select_out(sw_042_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_042_module_data_in[7] ,
    \sw_042_module_data_in[6] ,
    \sw_042_module_data_in[5] ,
    \sw_042_module_data_in[4] ,
    \sw_042_module_data_in[3] ,
    \sw_042_module_data_in[2] ,
    \sw_042_module_data_in[1] ,
    \sw_042_module_data_in[0] }),
    .module_data_out({\sw_042_module_data_out[7] ,
    \sw_042_module_data_out[6] ,
    \sw_042_module_data_out[5] ,
    \sw_042_module_data_out[4] ,
    \sw_042_module_data_out[3] ,
    \sw_042_module_data_out[2] ,
    \sw_042_module_data_out[1] ,
    \sw_042_module_data_out[0] }));
 scanchain scanchain_043 (.clk_in(sw_042_clk_out),
    .clk_out(sw_043_clk_out),
    .data_in(sw_042_data_out),
    .data_out(sw_043_data_out),
    .latch_enable_in(sw_042_latch_out),
    .latch_enable_out(sw_043_latch_out),
    .scan_select_in(sw_042_scan_out),
    .scan_select_out(sw_043_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_043_module_data_in[7] ,
    \sw_043_module_data_in[6] ,
    \sw_043_module_data_in[5] ,
    \sw_043_module_data_in[4] ,
    \sw_043_module_data_in[3] ,
    \sw_043_module_data_in[2] ,
    \sw_043_module_data_in[1] ,
    \sw_043_module_data_in[0] }),
    .module_data_out({\sw_043_module_data_out[7] ,
    \sw_043_module_data_out[6] ,
    \sw_043_module_data_out[5] ,
    \sw_043_module_data_out[4] ,
    \sw_043_module_data_out[3] ,
    \sw_043_module_data_out[2] ,
    \sw_043_module_data_out[1] ,
    \sw_043_module_data_out[0] }));
 scanchain scanchain_044 (.clk_in(sw_043_clk_out),
    .clk_out(sw_044_clk_out),
    .data_in(sw_043_data_out),
    .data_out(sw_044_data_out),
    .latch_enable_in(sw_043_latch_out),
    .latch_enable_out(sw_044_latch_out),
    .scan_select_in(sw_043_scan_out),
    .scan_select_out(sw_044_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_044_module_data_in[7] ,
    \sw_044_module_data_in[6] ,
    \sw_044_module_data_in[5] ,
    \sw_044_module_data_in[4] ,
    \sw_044_module_data_in[3] ,
    \sw_044_module_data_in[2] ,
    \sw_044_module_data_in[1] ,
    \sw_044_module_data_in[0] }),
    .module_data_out({\sw_044_module_data_out[7] ,
    \sw_044_module_data_out[6] ,
    \sw_044_module_data_out[5] ,
    \sw_044_module_data_out[4] ,
    \sw_044_module_data_out[3] ,
    \sw_044_module_data_out[2] ,
    \sw_044_module_data_out[1] ,
    \sw_044_module_data_out[0] }));
 scanchain scanchain_045 (.clk_in(sw_044_clk_out),
    .clk_out(sw_045_clk_out),
    .data_in(sw_044_data_out),
    .data_out(sw_045_data_out),
    .latch_enable_in(sw_044_latch_out),
    .latch_enable_out(sw_045_latch_out),
    .scan_select_in(sw_044_scan_out),
    .scan_select_out(sw_045_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_045_module_data_in[7] ,
    \sw_045_module_data_in[6] ,
    \sw_045_module_data_in[5] ,
    \sw_045_module_data_in[4] ,
    \sw_045_module_data_in[3] ,
    \sw_045_module_data_in[2] ,
    \sw_045_module_data_in[1] ,
    \sw_045_module_data_in[0] }),
    .module_data_out({\sw_045_module_data_out[7] ,
    \sw_045_module_data_out[6] ,
    \sw_045_module_data_out[5] ,
    \sw_045_module_data_out[4] ,
    \sw_045_module_data_out[3] ,
    \sw_045_module_data_out[2] ,
    \sw_045_module_data_out[1] ,
    \sw_045_module_data_out[0] }));
 scanchain scanchain_046 (.clk_in(sw_045_clk_out),
    .clk_out(sw_046_clk_out),
    .data_in(sw_045_data_out),
    .data_out(sw_046_data_out),
    .latch_enable_in(sw_045_latch_out),
    .latch_enable_out(sw_046_latch_out),
    .scan_select_in(sw_045_scan_out),
    .scan_select_out(sw_046_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_046_module_data_in[7] ,
    \sw_046_module_data_in[6] ,
    \sw_046_module_data_in[5] ,
    \sw_046_module_data_in[4] ,
    \sw_046_module_data_in[3] ,
    \sw_046_module_data_in[2] ,
    \sw_046_module_data_in[1] ,
    \sw_046_module_data_in[0] }),
    .module_data_out({\sw_046_module_data_out[7] ,
    \sw_046_module_data_out[6] ,
    \sw_046_module_data_out[5] ,
    \sw_046_module_data_out[4] ,
    \sw_046_module_data_out[3] ,
    \sw_046_module_data_out[2] ,
    \sw_046_module_data_out[1] ,
    \sw_046_module_data_out[0] }));
 scanchain scanchain_047 (.clk_in(sw_046_clk_out),
    .clk_out(sw_047_clk_out),
    .data_in(sw_046_data_out),
    .data_out(sw_047_data_out),
    .latch_enable_in(sw_046_latch_out),
    .latch_enable_out(sw_047_latch_out),
    .scan_select_in(sw_046_scan_out),
    .scan_select_out(sw_047_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_047_module_data_in[7] ,
    \sw_047_module_data_in[6] ,
    \sw_047_module_data_in[5] ,
    \sw_047_module_data_in[4] ,
    \sw_047_module_data_in[3] ,
    \sw_047_module_data_in[2] ,
    \sw_047_module_data_in[1] ,
    \sw_047_module_data_in[0] }),
    .module_data_out({\sw_047_module_data_out[7] ,
    \sw_047_module_data_out[6] ,
    \sw_047_module_data_out[5] ,
    \sw_047_module_data_out[4] ,
    \sw_047_module_data_out[3] ,
    \sw_047_module_data_out[2] ,
    \sw_047_module_data_out[1] ,
    \sw_047_module_data_out[0] }));
 scanchain scanchain_048 (.clk_in(sw_047_clk_out),
    .clk_out(sw_048_clk_out),
    .data_in(sw_047_data_out),
    .data_out(sw_048_data_out),
    .latch_enable_in(sw_047_latch_out),
    .latch_enable_out(sw_048_latch_out),
    .scan_select_in(sw_047_scan_out),
    .scan_select_out(sw_048_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_048_module_data_in[7] ,
    \sw_048_module_data_in[6] ,
    \sw_048_module_data_in[5] ,
    \sw_048_module_data_in[4] ,
    \sw_048_module_data_in[3] ,
    \sw_048_module_data_in[2] ,
    \sw_048_module_data_in[1] ,
    \sw_048_module_data_in[0] }),
    .module_data_out({\sw_048_module_data_out[7] ,
    \sw_048_module_data_out[6] ,
    \sw_048_module_data_out[5] ,
    \sw_048_module_data_out[4] ,
    \sw_048_module_data_out[3] ,
    \sw_048_module_data_out[2] ,
    \sw_048_module_data_out[1] ,
    \sw_048_module_data_out[0] }));
 scanchain scanchain_049 (.clk_in(sw_048_clk_out),
    .clk_out(sw_049_clk_out),
    .data_in(sw_048_data_out),
    .data_out(sw_049_data_out),
    .latch_enable_in(sw_048_latch_out),
    .latch_enable_out(sw_049_latch_out),
    .scan_select_in(sw_048_scan_out),
    .scan_select_out(sw_049_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_049_module_data_in[7] ,
    \sw_049_module_data_in[6] ,
    \sw_049_module_data_in[5] ,
    \sw_049_module_data_in[4] ,
    \sw_049_module_data_in[3] ,
    \sw_049_module_data_in[2] ,
    \sw_049_module_data_in[1] ,
    \sw_049_module_data_in[0] }),
    .module_data_out({\sw_049_module_data_out[7] ,
    \sw_049_module_data_out[6] ,
    \sw_049_module_data_out[5] ,
    \sw_049_module_data_out[4] ,
    \sw_049_module_data_out[3] ,
    \sw_049_module_data_out[2] ,
    \sw_049_module_data_out[1] ,
    \sw_049_module_data_out[0] }));
 scanchain scanchain_050 (.clk_in(sw_049_clk_out),
    .clk_out(sw_050_clk_out),
    .data_in(sw_049_data_out),
    .data_out(sw_050_data_out),
    .latch_enable_in(sw_049_latch_out),
    .latch_enable_out(sw_050_latch_out),
    .scan_select_in(sw_049_scan_out),
    .scan_select_out(sw_050_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_050_module_data_in[7] ,
    \sw_050_module_data_in[6] ,
    \sw_050_module_data_in[5] ,
    \sw_050_module_data_in[4] ,
    \sw_050_module_data_in[3] ,
    \sw_050_module_data_in[2] ,
    \sw_050_module_data_in[1] ,
    \sw_050_module_data_in[0] }),
    .module_data_out({\sw_050_module_data_out[7] ,
    \sw_050_module_data_out[6] ,
    \sw_050_module_data_out[5] ,
    \sw_050_module_data_out[4] ,
    \sw_050_module_data_out[3] ,
    \sw_050_module_data_out[2] ,
    \sw_050_module_data_out[1] ,
    \sw_050_module_data_out[0] }));
 scanchain scanchain_051 (.clk_in(sw_050_clk_out),
    .clk_out(sw_051_clk_out),
    .data_in(sw_050_data_out),
    .data_out(sw_051_data_out),
    .latch_enable_in(sw_050_latch_out),
    .latch_enable_out(sw_051_latch_out),
    .scan_select_in(sw_050_scan_out),
    .scan_select_out(sw_051_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_051_module_data_in[7] ,
    \sw_051_module_data_in[6] ,
    \sw_051_module_data_in[5] ,
    \sw_051_module_data_in[4] ,
    \sw_051_module_data_in[3] ,
    \sw_051_module_data_in[2] ,
    \sw_051_module_data_in[1] ,
    \sw_051_module_data_in[0] }),
    .module_data_out({\sw_051_module_data_out[7] ,
    \sw_051_module_data_out[6] ,
    \sw_051_module_data_out[5] ,
    \sw_051_module_data_out[4] ,
    \sw_051_module_data_out[3] ,
    \sw_051_module_data_out[2] ,
    \sw_051_module_data_out[1] ,
    \sw_051_module_data_out[0] }));
 scanchain scanchain_052 (.clk_in(sw_051_clk_out),
    .clk_out(sw_052_clk_out),
    .data_in(sw_051_data_out),
    .data_out(sw_052_data_out),
    .latch_enable_in(sw_051_latch_out),
    .latch_enable_out(sw_052_latch_out),
    .scan_select_in(sw_051_scan_out),
    .scan_select_out(sw_052_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_052_module_data_in[7] ,
    \sw_052_module_data_in[6] ,
    \sw_052_module_data_in[5] ,
    \sw_052_module_data_in[4] ,
    \sw_052_module_data_in[3] ,
    \sw_052_module_data_in[2] ,
    \sw_052_module_data_in[1] ,
    \sw_052_module_data_in[0] }),
    .module_data_out({\sw_052_module_data_out[7] ,
    \sw_052_module_data_out[6] ,
    \sw_052_module_data_out[5] ,
    \sw_052_module_data_out[4] ,
    \sw_052_module_data_out[3] ,
    \sw_052_module_data_out[2] ,
    \sw_052_module_data_out[1] ,
    \sw_052_module_data_out[0] }));
 scanchain scanchain_053 (.clk_in(sw_052_clk_out),
    .clk_out(sw_053_clk_out),
    .data_in(sw_052_data_out),
    .data_out(sw_053_data_out),
    .latch_enable_in(sw_052_latch_out),
    .latch_enable_out(sw_053_latch_out),
    .scan_select_in(sw_052_scan_out),
    .scan_select_out(sw_053_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_053_module_data_in[7] ,
    \sw_053_module_data_in[6] ,
    \sw_053_module_data_in[5] ,
    \sw_053_module_data_in[4] ,
    \sw_053_module_data_in[3] ,
    \sw_053_module_data_in[2] ,
    \sw_053_module_data_in[1] ,
    \sw_053_module_data_in[0] }),
    .module_data_out({\sw_053_module_data_out[7] ,
    \sw_053_module_data_out[6] ,
    \sw_053_module_data_out[5] ,
    \sw_053_module_data_out[4] ,
    \sw_053_module_data_out[3] ,
    \sw_053_module_data_out[2] ,
    \sw_053_module_data_out[1] ,
    \sw_053_module_data_out[0] }));
 scanchain scanchain_054 (.clk_in(sw_053_clk_out),
    .clk_out(sw_054_clk_out),
    .data_in(sw_053_data_out),
    .data_out(sw_054_data_out),
    .latch_enable_in(sw_053_latch_out),
    .latch_enable_out(sw_054_latch_out),
    .scan_select_in(sw_053_scan_out),
    .scan_select_out(sw_054_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_054_module_data_in[7] ,
    \sw_054_module_data_in[6] ,
    \sw_054_module_data_in[5] ,
    \sw_054_module_data_in[4] ,
    \sw_054_module_data_in[3] ,
    \sw_054_module_data_in[2] ,
    \sw_054_module_data_in[1] ,
    \sw_054_module_data_in[0] }),
    .module_data_out({\sw_054_module_data_out[7] ,
    \sw_054_module_data_out[6] ,
    \sw_054_module_data_out[5] ,
    \sw_054_module_data_out[4] ,
    \sw_054_module_data_out[3] ,
    \sw_054_module_data_out[2] ,
    \sw_054_module_data_out[1] ,
    \sw_054_module_data_out[0] }));
 scanchain scanchain_055 (.clk_in(sw_054_clk_out),
    .clk_out(sw_055_clk_out),
    .data_in(sw_054_data_out),
    .data_out(sw_055_data_out),
    .latch_enable_in(sw_054_latch_out),
    .latch_enable_out(sw_055_latch_out),
    .scan_select_in(sw_054_scan_out),
    .scan_select_out(sw_055_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_055_module_data_in[7] ,
    \sw_055_module_data_in[6] ,
    \sw_055_module_data_in[5] ,
    \sw_055_module_data_in[4] ,
    \sw_055_module_data_in[3] ,
    \sw_055_module_data_in[2] ,
    \sw_055_module_data_in[1] ,
    \sw_055_module_data_in[0] }),
    .module_data_out({\sw_055_module_data_out[7] ,
    \sw_055_module_data_out[6] ,
    \sw_055_module_data_out[5] ,
    \sw_055_module_data_out[4] ,
    \sw_055_module_data_out[3] ,
    \sw_055_module_data_out[2] ,
    \sw_055_module_data_out[1] ,
    \sw_055_module_data_out[0] }));
 scanchain scanchain_056 (.clk_in(sw_055_clk_out),
    .clk_out(sw_056_clk_out),
    .data_in(sw_055_data_out),
    .data_out(sw_056_data_out),
    .latch_enable_in(sw_055_latch_out),
    .latch_enable_out(sw_056_latch_out),
    .scan_select_in(sw_055_scan_out),
    .scan_select_out(sw_056_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_056_module_data_in[7] ,
    \sw_056_module_data_in[6] ,
    \sw_056_module_data_in[5] ,
    \sw_056_module_data_in[4] ,
    \sw_056_module_data_in[3] ,
    \sw_056_module_data_in[2] ,
    \sw_056_module_data_in[1] ,
    \sw_056_module_data_in[0] }),
    .module_data_out({\sw_056_module_data_out[7] ,
    \sw_056_module_data_out[6] ,
    \sw_056_module_data_out[5] ,
    \sw_056_module_data_out[4] ,
    \sw_056_module_data_out[3] ,
    \sw_056_module_data_out[2] ,
    \sw_056_module_data_out[1] ,
    \sw_056_module_data_out[0] }));
 scanchain scanchain_057 (.clk_in(sw_056_clk_out),
    .clk_out(sw_057_clk_out),
    .data_in(sw_056_data_out),
    .data_out(sw_057_data_out),
    .latch_enable_in(sw_056_latch_out),
    .latch_enable_out(sw_057_latch_out),
    .scan_select_in(sw_056_scan_out),
    .scan_select_out(sw_057_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_057_module_data_in[7] ,
    \sw_057_module_data_in[6] ,
    \sw_057_module_data_in[5] ,
    \sw_057_module_data_in[4] ,
    \sw_057_module_data_in[3] ,
    \sw_057_module_data_in[2] ,
    \sw_057_module_data_in[1] ,
    \sw_057_module_data_in[0] }),
    .module_data_out({\sw_057_module_data_out[7] ,
    \sw_057_module_data_out[6] ,
    \sw_057_module_data_out[5] ,
    \sw_057_module_data_out[4] ,
    \sw_057_module_data_out[3] ,
    \sw_057_module_data_out[2] ,
    \sw_057_module_data_out[1] ,
    \sw_057_module_data_out[0] }));
 scanchain scanchain_058 (.clk_in(sw_057_clk_out),
    .clk_out(sw_058_clk_out),
    .data_in(sw_057_data_out),
    .data_out(sw_058_data_out),
    .latch_enable_in(sw_057_latch_out),
    .latch_enable_out(sw_058_latch_out),
    .scan_select_in(sw_057_scan_out),
    .scan_select_out(sw_058_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_058_module_data_in[7] ,
    \sw_058_module_data_in[6] ,
    \sw_058_module_data_in[5] ,
    \sw_058_module_data_in[4] ,
    \sw_058_module_data_in[3] ,
    \sw_058_module_data_in[2] ,
    \sw_058_module_data_in[1] ,
    \sw_058_module_data_in[0] }),
    .module_data_out({\sw_058_module_data_out[7] ,
    \sw_058_module_data_out[6] ,
    \sw_058_module_data_out[5] ,
    \sw_058_module_data_out[4] ,
    \sw_058_module_data_out[3] ,
    \sw_058_module_data_out[2] ,
    \sw_058_module_data_out[1] ,
    \sw_058_module_data_out[0] }));
 scanchain scanchain_059 (.clk_in(sw_058_clk_out),
    .clk_out(sw_059_clk_out),
    .data_in(sw_058_data_out),
    .data_out(sw_059_data_out),
    .latch_enable_in(sw_058_latch_out),
    .latch_enable_out(sw_059_latch_out),
    .scan_select_in(sw_058_scan_out),
    .scan_select_out(sw_059_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_059_module_data_in[7] ,
    \sw_059_module_data_in[6] ,
    \sw_059_module_data_in[5] ,
    \sw_059_module_data_in[4] ,
    \sw_059_module_data_in[3] ,
    \sw_059_module_data_in[2] ,
    \sw_059_module_data_in[1] ,
    \sw_059_module_data_in[0] }),
    .module_data_out({\sw_059_module_data_out[7] ,
    \sw_059_module_data_out[6] ,
    \sw_059_module_data_out[5] ,
    \sw_059_module_data_out[4] ,
    \sw_059_module_data_out[3] ,
    \sw_059_module_data_out[2] ,
    \sw_059_module_data_out[1] ,
    \sw_059_module_data_out[0] }));
 scanchain scanchain_060 (.clk_in(sw_059_clk_out),
    .clk_out(sw_060_clk_out),
    .data_in(sw_059_data_out),
    .data_out(sw_060_data_out),
    .latch_enable_in(sw_059_latch_out),
    .latch_enable_out(sw_060_latch_out),
    .scan_select_in(sw_059_scan_out),
    .scan_select_out(sw_060_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_060_module_data_in[7] ,
    \sw_060_module_data_in[6] ,
    \sw_060_module_data_in[5] ,
    \sw_060_module_data_in[4] ,
    \sw_060_module_data_in[3] ,
    \sw_060_module_data_in[2] ,
    \sw_060_module_data_in[1] ,
    \sw_060_module_data_in[0] }),
    .module_data_out({\sw_060_module_data_out[7] ,
    \sw_060_module_data_out[6] ,
    \sw_060_module_data_out[5] ,
    \sw_060_module_data_out[4] ,
    \sw_060_module_data_out[3] ,
    \sw_060_module_data_out[2] ,
    \sw_060_module_data_out[1] ,
    \sw_060_module_data_out[0] }));
 scanchain scanchain_061 (.clk_in(sw_060_clk_out),
    .clk_out(sw_061_clk_out),
    .data_in(sw_060_data_out),
    .data_out(sw_061_data_out),
    .latch_enable_in(sw_060_latch_out),
    .latch_enable_out(sw_061_latch_out),
    .scan_select_in(sw_060_scan_out),
    .scan_select_out(sw_061_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_061_module_data_in[7] ,
    \sw_061_module_data_in[6] ,
    \sw_061_module_data_in[5] ,
    \sw_061_module_data_in[4] ,
    \sw_061_module_data_in[3] ,
    \sw_061_module_data_in[2] ,
    \sw_061_module_data_in[1] ,
    \sw_061_module_data_in[0] }),
    .module_data_out({\sw_061_module_data_out[7] ,
    \sw_061_module_data_out[6] ,
    \sw_061_module_data_out[5] ,
    \sw_061_module_data_out[4] ,
    \sw_061_module_data_out[3] ,
    \sw_061_module_data_out[2] ,
    \sw_061_module_data_out[1] ,
    \sw_061_module_data_out[0] }));
 scanchain scanchain_062 (.clk_in(sw_061_clk_out),
    .clk_out(sw_062_clk_out),
    .data_in(sw_061_data_out),
    .data_out(sw_062_data_out),
    .latch_enable_in(sw_061_latch_out),
    .latch_enable_out(sw_062_latch_out),
    .scan_select_in(sw_061_scan_out),
    .scan_select_out(sw_062_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_062_module_data_in[7] ,
    \sw_062_module_data_in[6] ,
    \sw_062_module_data_in[5] ,
    \sw_062_module_data_in[4] ,
    \sw_062_module_data_in[3] ,
    \sw_062_module_data_in[2] ,
    \sw_062_module_data_in[1] ,
    \sw_062_module_data_in[0] }),
    .module_data_out({\sw_062_module_data_out[7] ,
    \sw_062_module_data_out[6] ,
    \sw_062_module_data_out[5] ,
    \sw_062_module_data_out[4] ,
    \sw_062_module_data_out[3] ,
    \sw_062_module_data_out[2] ,
    \sw_062_module_data_out[1] ,
    \sw_062_module_data_out[0] }));
 scanchain scanchain_063 (.clk_in(sw_062_clk_out),
    .clk_out(sw_063_clk_out),
    .data_in(sw_062_data_out),
    .data_out(sw_063_data_out),
    .latch_enable_in(sw_062_latch_out),
    .latch_enable_out(sw_063_latch_out),
    .scan_select_in(sw_062_scan_out),
    .scan_select_out(sw_063_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_063_module_data_in[7] ,
    \sw_063_module_data_in[6] ,
    \sw_063_module_data_in[5] ,
    \sw_063_module_data_in[4] ,
    \sw_063_module_data_in[3] ,
    \sw_063_module_data_in[2] ,
    \sw_063_module_data_in[1] ,
    \sw_063_module_data_in[0] }),
    .module_data_out({\sw_063_module_data_out[7] ,
    \sw_063_module_data_out[6] ,
    \sw_063_module_data_out[5] ,
    \sw_063_module_data_out[4] ,
    \sw_063_module_data_out[3] ,
    \sw_063_module_data_out[2] ,
    \sw_063_module_data_out[1] ,
    \sw_063_module_data_out[0] }));
 scanchain scanchain_064 (.clk_in(sw_063_clk_out),
    .clk_out(sw_064_clk_out),
    .data_in(sw_063_data_out),
    .data_out(sw_064_data_out),
    .latch_enable_in(sw_063_latch_out),
    .latch_enable_out(sw_064_latch_out),
    .scan_select_in(sw_063_scan_out),
    .scan_select_out(sw_064_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_064_module_data_in[7] ,
    \sw_064_module_data_in[6] ,
    \sw_064_module_data_in[5] ,
    \sw_064_module_data_in[4] ,
    \sw_064_module_data_in[3] ,
    \sw_064_module_data_in[2] ,
    \sw_064_module_data_in[1] ,
    \sw_064_module_data_in[0] }),
    .module_data_out({\sw_064_module_data_out[7] ,
    \sw_064_module_data_out[6] ,
    \sw_064_module_data_out[5] ,
    \sw_064_module_data_out[4] ,
    \sw_064_module_data_out[3] ,
    \sw_064_module_data_out[2] ,
    \sw_064_module_data_out[1] ,
    \sw_064_module_data_out[0] }));
 scanchain scanchain_065 (.clk_in(sw_064_clk_out),
    .clk_out(sw_065_clk_out),
    .data_in(sw_064_data_out),
    .data_out(sw_065_data_out),
    .latch_enable_in(sw_064_latch_out),
    .latch_enable_out(sw_065_latch_out),
    .scan_select_in(sw_064_scan_out),
    .scan_select_out(sw_065_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_065_module_data_in[7] ,
    \sw_065_module_data_in[6] ,
    \sw_065_module_data_in[5] ,
    \sw_065_module_data_in[4] ,
    \sw_065_module_data_in[3] ,
    \sw_065_module_data_in[2] ,
    \sw_065_module_data_in[1] ,
    \sw_065_module_data_in[0] }),
    .module_data_out({\sw_065_module_data_out[7] ,
    \sw_065_module_data_out[6] ,
    \sw_065_module_data_out[5] ,
    \sw_065_module_data_out[4] ,
    \sw_065_module_data_out[3] ,
    \sw_065_module_data_out[2] ,
    \sw_065_module_data_out[1] ,
    \sw_065_module_data_out[0] }));
 scanchain scanchain_066 (.clk_in(sw_065_clk_out),
    .clk_out(sw_066_clk_out),
    .data_in(sw_065_data_out),
    .data_out(sw_066_data_out),
    .latch_enable_in(sw_065_latch_out),
    .latch_enable_out(sw_066_latch_out),
    .scan_select_in(sw_065_scan_out),
    .scan_select_out(sw_066_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_066_module_data_in[7] ,
    \sw_066_module_data_in[6] ,
    \sw_066_module_data_in[5] ,
    \sw_066_module_data_in[4] ,
    \sw_066_module_data_in[3] ,
    \sw_066_module_data_in[2] ,
    \sw_066_module_data_in[1] ,
    \sw_066_module_data_in[0] }),
    .module_data_out({\sw_066_module_data_out[7] ,
    \sw_066_module_data_out[6] ,
    \sw_066_module_data_out[5] ,
    \sw_066_module_data_out[4] ,
    \sw_066_module_data_out[3] ,
    \sw_066_module_data_out[2] ,
    \sw_066_module_data_out[1] ,
    \sw_066_module_data_out[0] }));
 scanchain scanchain_067 (.clk_in(sw_066_clk_out),
    .clk_out(sw_067_clk_out),
    .data_in(sw_066_data_out),
    .data_out(sw_067_data_out),
    .latch_enable_in(sw_066_latch_out),
    .latch_enable_out(sw_067_latch_out),
    .scan_select_in(sw_066_scan_out),
    .scan_select_out(sw_067_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_067_module_data_in[7] ,
    \sw_067_module_data_in[6] ,
    \sw_067_module_data_in[5] ,
    \sw_067_module_data_in[4] ,
    \sw_067_module_data_in[3] ,
    \sw_067_module_data_in[2] ,
    \sw_067_module_data_in[1] ,
    \sw_067_module_data_in[0] }),
    .module_data_out({\sw_067_module_data_out[7] ,
    \sw_067_module_data_out[6] ,
    \sw_067_module_data_out[5] ,
    \sw_067_module_data_out[4] ,
    \sw_067_module_data_out[3] ,
    \sw_067_module_data_out[2] ,
    \sw_067_module_data_out[1] ,
    \sw_067_module_data_out[0] }));
 scanchain scanchain_068 (.clk_in(sw_067_clk_out),
    .clk_out(sw_068_clk_out),
    .data_in(sw_067_data_out),
    .data_out(sw_068_data_out),
    .latch_enable_in(sw_067_latch_out),
    .latch_enable_out(sw_068_latch_out),
    .scan_select_in(sw_067_scan_out),
    .scan_select_out(sw_068_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_068_module_data_in[7] ,
    \sw_068_module_data_in[6] ,
    \sw_068_module_data_in[5] ,
    \sw_068_module_data_in[4] ,
    \sw_068_module_data_in[3] ,
    \sw_068_module_data_in[2] ,
    \sw_068_module_data_in[1] ,
    \sw_068_module_data_in[0] }),
    .module_data_out({\sw_068_module_data_out[7] ,
    \sw_068_module_data_out[6] ,
    \sw_068_module_data_out[5] ,
    \sw_068_module_data_out[4] ,
    \sw_068_module_data_out[3] ,
    \sw_068_module_data_out[2] ,
    \sw_068_module_data_out[1] ,
    \sw_068_module_data_out[0] }));
 scanchain scanchain_069 (.clk_in(sw_068_clk_out),
    .clk_out(sw_069_clk_out),
    .data_in(sw_068_data_out),
    .data_out(sw_069_data_out),
    .latch_enable_in(sw_068_latch_out),
    .latch_enable_out(sw_069_latch_out),
    .scan_select_in(sw_068_scan_out),
    .scan_select_out(sw_069_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_069_module_data_in[7] ,
    \sw_069_module_data_in[6] ,
    \sw_069_module_data_in[5] ,
    \sw_069_module_data_in[4] ,
    \sw_069_module_data_in[3] ,
    \sw_069_module_data_in[2] ,
    \sw_069_module_data_in[1] ,
    \sw_069_module_data_in[0] }),
    .module_data_out({\sw_069_module_data_out[7] ,
    \sw_069_module_data_out[6] ,
    \sw_069_module_data_out[5] ,
    \sw_069_module_data_out[4] ,
    \sw_069_module_data_out[3] ,
    \sw_069_module_data_out[2] ,
    \sw_069_module_data_out[1] ,
    \sw_069_module_data_out[0] }));
 scanchain scanchain_070 (.clk_in(sw_069_clk_out),
    .clk_out(sw_070_clk_out),
    .data_in(sw_069_data_out),
    .data_out(sw_070_data_out),
    .latch_enable_in(sw_069_latch_out),
    .latch_enable_out(sw_070_latch_out),
    .scan_select_in(sw_069_scan_out),
    .scan_select_out(sw_070_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_070_module_data_in[7] ,
    \sw_070_module_data_in[6] ,
    \sw_070_module_data_in[5] ,
    \sw_070_module_data_in[4] ,
    \sw_070_module_data_in[3] ,
    \sw_070_module_data_in[2] ,
    \sw_070_module_data_in[1] ,
    \sw_070_module_data_in[0] }),
    .module_data_out({\sw_070_module_data_out[7] ,
    \sw_070_module_data_out[6] ,
    \sw_070_module_data_out[5] ,
    \sw_070_module_data_out[4] ,
    \sw_070_module_data_out[3] ,
    \sw_070_module_data_out[2] ,
    \sw_070_module_data_out[1] ,
    \sw_070_module_data_out[0] }));
 scanchain scanchain_071 (.clk_in(sw_070_clk_out),
    .clk_out(sw_071_clk_out),
    .data_in(sw_070_data_out),
    .data_out(sw_071_data_out),
    .latch_enable_in(sw_070_latch_out),
    .latch_enable_out(sw_071_latch_out),
    .scan_select_in(sw_070_scan_out),
    .scan_select_out(sw_071_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_071_module_data_in[7] ,
    \sw_071_module_data_in[6] ,
    \sw_071_module_data_in[5] ,
    \sw_071_module_data_in[4] ,
    \sw_071_module_data_in[3] ,
    \sw_071_module_data_in[2] ,
    \sw_071_module_data_in[1] ,
    \sw_071_module_data_in[0] }),
    .module_data_out({\sw_071_module_data_out[7] ,
    \sw_071_module_data_out[6] ,
    \sw_071_module_data_out[5] ,
    \sw_071_module_data_out[4] ,
    \sw_071_module_data_out[3] ,
    \sw_071_module_data_out[2] ,
    \sw_071_module_data_out[1] ,
    \sw_071_module_data_out[0] }));
 scanchain scanchain_072 (.clk_in(sw_071_clk_out),
    .clk_out(sw_072_clk_out),
    .data_in(sw_071_data_out),
    .data_out(sw_072_data_out),
    .latch_enable_in(sw_071_latch_out),
    .latch_enable_out(sw_072_latch_out),
    .scan_select_in(sw_071_scan_out),
    .scan_select_out(sw_072_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_072_module_data_in[7] ,
    \sw_072_module_data_in[6] ,
    \sw_072_module_data_in[5] ,
    \sw_072_module_data_in[4] ,
    \sw_072_module_data_in[3] ,
    \sw_072_module_data_in[2] ,
    \sw_072_module_data_in[1] ,
    \sw_072_module_data_in[0] }),
    .module_data_out({\sw_072_module_data_out[7] ,
    \sw_072_module_data_out[6] ,
    \sw_072_module_data_out[5] ,
    \sw_072_module_data_out[4] ,
    \sw_072_module_data_out[3] ,
    \sw_072_module_data_out[2] ,
    \sw_072_module_data_out[1] ,
    \sw_072_module_data_out[0] }));
 scanchain scanchain_073 (.clk_in(sw_072_clk_out),
    .clk_out(sw_073_clk_out),
    .data_in(sw_072_data_out),
    .data_out(sw_073_data_out),
    .latch_enable_in(sw_072_latch_out),
    .latch_enable_out(sw_073_latch_out),
    .scan_select_in(sw_072_scan_out),
    .scan_select_out(sw_073_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_073_module_data_in[7] ,
    \sw_073_module_data_in[6] ,
    \sw_073_module_data_in[5] ,
    \sw_073_module_data_in[4] ,
    \sw_073_module_data_in[3] ,
    \sw_073_module_data_in[2] ,
    \sw_073_module_data_in[1] ,
    \sw_073_module_data_in[0] }),
    .module_data_out({\sw_073_module_data_out[7] ,
    \sw_073_module_data_out[6] ,
    \sw_073_module_data_out[5] ,
    \sw_073_module_data_out[4] ,
    \sw_073_module_data_out[3] ,
    \sw_073_module_data_out[2] ,
    \sw_073_module_data_out[1] ,
    \sw_073_module_data_out[0] }));
 scanchain scanchain_074 (.clk_in(sw_073_clk_out),
    .clk_out(sw_074_clk_out),
    .data_in(sw_073_data_out),
    .data_out(sw_074_data_out),
    .latch_enable_in(sw_073_latch_out),
    .latch_enable_out(sw_074_latch_out),
    .scan_select_in(sw_073_scan_out),
    .scan_select_out(sw_074_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_074_module_data_in[7] ,
    \sw_074_module_data_in[6] ,
    \sw_074_module_data_in[5] ,
    \sw_074_module_data_in[4] ,
    \sw_074_module_data_in[3] ,
    \sw_074_module_data_in[2] ,
    \sw_074_module_data_in[1] ,
    \sw_074_module_data_in[0] }),
    .module_data_out({\sw_074_module_data_out[7] ,
    \sw_074_module_data_out[6] ,
    \sw_074_module_data_out[5] ,
    \sw_074_module_data_out[4] ,
    \sw_074_module_data_out[3] ,
    \sw_074_module_data_out[2] ,
    \sw_074_module_data_out[1] ,
    \sw_074_module_data_out[0] }));
 scanchain scanchain_075 (.clk_in(sw_074_clk_out),
    .clk_out(sw_075_clk_out),
    .data_in(sw_074_data_out),
    .data_out(sw_075_data_out),
    .latch_enable_in(sw_074_latch_out),
    .latch_enable_out(sw_075_latch_out),
    .scan_select_in(sw_074_scan_out),
    .scan_select_out(sw_075_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_075_module_data_in[7] ,
    \sw_075_module_data_in[6] ,
    \sw_075_module_data_in[5] ,
    \sw_075_module_data_in[4] ,
    \sw_075_module_data_in[3] ,
    \sw_075_module_data_in[2] ,
    \sw_075_module_data_in[1] ,
    \sw_075_module_data_in[0] }),
    .module_data_out({\sw_075_module_data_out[7] ,
    \sw_075_module_data_out[6] ,
    \sw_075_module_data_out[5] ,
    \sw_075_module_data_out[4] ,
    \sw_075_module_data_out[3] ,
    \sw_075_module_data_out[2] ,
    \sw_075_module_data_out[1] ,
    \sw_075_module_data_out[0] }));
 scanchain scanchain_076 (.clk_in(sw_075_clk_out),
    .clk_out(sw_076_clk_out),
    .data_in(sw_075_data_out),
    .data_out(sw_076_data_out),
    .latch_enable_in(sw_075_latch_out),
    .latch_enable_out(sw_076_latch_out),
    .scan_select_in(sw_075_scan_out),
    .scan_select_out(sw_076_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_076_module_data_in[7] ,
    \sw_076_module_data_in[6] ,
    \sw_076_module_data_in[5] ,
    \sw_076_module_data_in[4] ,
    \sw_076_module_data_in[3] ,
    \sw_076_module_data_in[2] ,
    \sw_076_module_data_in[1] ,
    \sw_076_module_data_in[0] }),
    .module_data_out({\sw_076_module_data_out[7] ,
    \sw_076_module_data_out[6] ,
    \sw_076_module_data_out[5] ,
    \sw_076_module_data_out[4] ,
    \sw_076_module_data_out[3] ,
    \sw_076_module_data_out[2] ,
    \sw_076_module_data_out[1] ,
    \sw_076_module_data_out[0] }));
 scanchain scanchain_077 (.clk_in(sw_076_clk_out),
    .clk_out(sw_077_clk_out),
    .data_in(sw_076_data_out),
    .data_out(sw_077_data_out),
    .latch_enable_in(sw_076_latch_out),
    .latch_enable_out(sw_077_latch_out),
    .scan_select_in(sw_076_scan_out),
    .scan_select_out(sw_077_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_077_module_data_in[7] ,
    \sw_077_module_data_in[6] ,
    \sw_077_module_data_in[5] ,
    \sw_077_module_data_in[4] ,
    \sw_077_module_data_in[3] ,
    \sw_077_module_data_in[2] ,
    \sw_077_module_data_in[1] ,
    \sw_077_module_data_in[0] }),
    .module_data_out({\sw_077_module_data_out[7] ,
    \sw_077_module_data_out[6] ,
    \sw_077_module_data_out[5] ,
    \sw_077_module_data_out[4] ,
    \sw_077_module_data_out[3] ,
    \sw_077_module_data_out[2] ,
    \sw_077_module_data_out[1] ,
    \sw_077_module_data_out[0] }));
 scanchain scanchain_078 (.clk_in(sw_077_clk_out),
    .clk_out(sw_078_clk_out),
    .data_in(sw_077_data_out),
    .data_out(sw_078_data_out),
    .latch_enable_in(sw_077_latch_out),
    .latch_enable_out(sw_078_latch_out),
    .scan_select_in(sw_077_scan_out),
    .scan_select_out(sw_078_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_078_module_data_in[7] ,
    \sw_078_module_data_in[6] ,
    \sw_078_module_data_in[5] ,
    \sw_078_module_data_in[4] ,
    \sw_078_module_data_in[3] ,
    \sw_078_module_data_in[2] ,
    \sw_078_module_data_in[1] ,
    \sw_078_module_data_in[0] }),
    .module_data_out({\sw_078_module_data_out[7] ,
    \sw_078_module_data_out[6] ,
    \sw_078_module_data_out[5] ,
    \sw_078_module_data_out[4] ,
    \sw_078_module_data_out[3] ,
    \sw_078_module_data_out[2] ,
    \sw_078_module_data_out[1] ,
    \sw_078_module_data_out[0] }));
 scanchain scanchain_079 (.clk_in(sw_078_clk_out),
    .clk_out(sw_079_clk_out),
    .data_in(sw_078_data_out),
    .data_out(sw_079_data_out),
    .latch_enable_in(sw_078_latch_out),
    .latch_enable_out(sw_079_latch_out),
    .scan_select_in(sw_078_scan_out),
    .scan_select_out(sw_079_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_079_module_data_in[7] ,
    \sw_079_module_data_in[6] ,
    \sw_079_module_data_in[5] ,
    \sw_079_module_data_in[4] ,
    \sw_079_module_data_in[3] ,
    \sw_079_module_data_in[2] ,
    \sw_079_module_data_in[1] ,
    \sw_079_module_data_in[0] }),
    .module_data_out({\sw_079_module_data_out[7] ,
    \sw_079_module_data_out[6] ,
    \sw_079_module_data_out[5] ,
    \sw_079_module_data_out[4] ,
    \sw_079_module_data_out[3] ,
    \sw_079_module_data_out[2] ,
    \sw_079_module_data_out[1] ,
    \sw_079_module_data_out[0] }));
 scanchain scanchain_080 (.clk_in(sw_079_clk_out),
    .clk_out(sw_080_clk_out),
    .data_in(sw_079_data_out),
    .data_out(sw_080_data_out),
    .latch_enable_in(sw_079_latch_out),
    .latch_enable_out(sw_080_latch_out),
    .scan_select_in(sw_079_scan_out),
    .scan_select_out(sw_080_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_080_module_data_in[7] ,
    \sw_080_module_data_in[6] ,
    \sw_080_module_data_in[5] ,
    \sw_080_module_data_in[4] ,
    \sw_080_module_data_in[3] ,
    \sw_080_module_data_in[2] ,
    \sw_080_module_data_in[1] ,
    \sw_080_module_data_in[0] }),
    .module_data_out({\sw_080_module_data_out[7] ,
    \sw_080_module_data_out[6] ,
    \sw_080_module_data_out[5] ,
    \sw_080_module_data_out[4] ,
    \sw_080_module_data_out[3] ,
    \sw_080_module_data_out[2] ,
    \sw_080_module_data_out[1] ,
    \sw_080_module_data_out[0] }));
 scanchain scanchain_081 (.clk_in(sw_080_clk_out),
    .clk_out(sw_081_clk_out),
    .data_in(sw_080_data_out),
    .data_out(sw_081_data_out),
    .latch_enable_in(sw_080_latch_out),
    .latch_enable_out(sw_081_latch_out),
    .scan_select_in(sw_080_scan_out),
    .scan_select_out(sw_081_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_081_module_data_in[7] ,
    \sw_081_module_data_in[6] ,
    \sw_081_module_data_in[5] ,
    \sw_081_module_data_in[4] ,
    \sw_081_module_data_in[3] ,
    \sw_081_module_data_in[2] ,
    \sw_081_module_data_in[1] ,
    \sw_081_module_data_in[0] }),
    .module_data_out({\sw_081_module_data_out[7] ,
    \sw_081_module_data_out[6] ,
    \sw_081_module_data_out[5] ,
    \sw_081_module_data_out[4] ,
    \sw_081_module_data_out[3] ,
    \sw_081_module_data_out[2] ,
    \sw_081_module_data_out[1] ,
    \sw_081_module_data_out[0] }));
 scanchain scanchain_082 (.clk_in(sw_081_clk_out),
    .clk_out(sw_082_clk_out),
    .data_in(sw_081_data_out),
    .data_out(sw_082_data_out),
    .latch_enable_in(sw_081_latch_out),
    .latch_enable_out(sw_082_latch_out),
    .scan_select_in(sw_081_scan_out),
    .scan_select_out(sw_082_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_082_module_data_in[7] ,
    \sw_082_module_data_in[6] ,
    \sw_082_module_data_in[5] ,
    \sw_082_module_data_in[4] ,
    \sw_082_module_data_in[3] ,
    \sw_082_module_data_in[2] ,
    \sw_082_module_data_in[1] ,
    \sw_082_module_data_in[0] }),
    .module_data_out({\sw_082_module_data_out[7] ,
    \sw_082_module_data_out[6] ,
    \sw_082_module_data_out[5] ,
    \sw_082_module_data_out[4] ,
    \sw_082_module_data_out[3] ,
    \sw_082_module_data_out[2] ,
    \sw_082_module_data_out[1] ,
    \sw_082_module_data_out[0] }));
 scanchain scanchain_083 (.clk_in(sw_082_clk_out),
    .clk_out(sw_083_clk_out),
    .data_in(sw_082_data_out),
    .data_out(sw_083_data_out),
    .latch_enable_in(sw_082_latch_out),
    .latch_enable_out(sw_083_latch_out),
    .scan_select_in(sw_082_scan_out),
    .scan_select_out(sw_083_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_083_module_data_in[7] ,
    \sw_083_module_data_in[6] ,
    \sw_083_module_data_in[5] ,
    \sw_083_module_data_in[4] ,
    \sw_083_module_data_in[3] ,
    \sw_083_module_data_in[2] ,
    \sw_083_module_data_in[1] ,
    \sw_083_module_data_in[0] }),
    .module_data_out({\sw_083_module_data_out[7] ,
    \sw_083_module_data_out[6] ,
    \sw_083_module_data_out[5] ,
    \sw_083_module_data_out[4] ,
    \sw_083_module_data_out[3] ,
    \sw_083_module_data_out[2] ,
    \sw_083_module_data_out[1] ,
    \sw_083_module_data_out[0] }));
 scanchain scanchain_084 (.clk_in(sw_083_clk_out),
    .clk_out(sw_084_clk_out),
    .data_in(sw_083_data_out),
    .data_out(sw_084_data_out),
    .latch_enable_in(sw_083_latch_out),
    .latch_enable_out(sw_084_latch_out),
    .scan_select_in(sw_083_scan_out),
    .scan_select_out(sw_084_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_084_module_data_in[7] ,
    \sw_084_module_data_in[6] ,
    \sw_084_module_data_in[5] ,
    \sw_084_module_data_in[4] ,
    \sw_084_module_data_in[3] ,
    \sw_084_module_data_in[2] ,
    \sw_084_module_data_in[1] ,
    \sw_084_module_data_in[0] }),
    .module_data_out({\sw_084_module_data_out[7] ,
    \sw_084_module_data_out[6] ,
    \sw_084_module_data_out[5] ,
    \sw_084_module_data_out[4] ,
    \sw_084_module_data_out[3] ,
    \sw_084_module_data_out[2] ,
    \sw_084_module_data_out[1] ,
    \sw_084_module_data_out[0] }));
 scanchain scanchain_085 (.clk_in(sw_084_clk_out),
    .clk_out(sw_085_clk_out),
    .data_in(sw_084_data_out),
    .data_out(sw_085_data_out),
    .latch_enable_in(sw_084_latch_out),
    .latch_enable_out(sw_085_latch_out),
    .scan_select_in(sw_084_scan_out),
    .scan_select_out(sw_085_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_085_module_data_in[7] ,
    \sw_085_module_data_in[6] ,
    \sw_085_module_data_in[5] ,
    \sw_085_module_data_in[4] ,
    \sw_085_module_data_in[3] ,
    \sw_085_module_data_in[2] ,
    \sw_085_module_data_in[1] ,
    \sw_085_module_data_in[0] }),
    .module_data_out({\sw_085_module_data_out[7] ,
    \sw_085_module_data_out[6] ,
    \sw_085_module_data_out[5] ,
    \sw_085_module_data_out[4] ,
    \sw_085_module_data_out[3] ,
    \sw_085_module_data_out[2] ,
    \sw_085_module_data_out[1] ,
    \sw_085_module_data_out[0] }));
 scanchain scanchain_086 (.clk_in(sw_085_clk_out),
    .clk_out(sw_086_clk_out),
    .data_in(sw_085_data_out),
    .data_out(sw_086_data_out),
    .latch_enable_in(sw_085_latch_out),
    .latch_enable_out(sw_086_latch_out),
    .scan_select_in(sw_085_scan_out),
    .scan_select_out(sw_086_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_086_module_data_in[7] ,
    \sw_086_module_data_in[6] ,
    \sw_086_module_data_in[5] ,
    \sw_086_module_data_in[4] ,
    \sw_086_module_data_in[3] ,
    \sw_086_module_data_in[2] ,
    \sw_086_module_data_in[1] ,
    \sw_086_module_data_in[0] }),
    .module_data_out({\sw_086_module_data_out[7] ,
    \sw_086_module_data_out[6] ,
    \sw_086_module_data_out[5] ,
    \sw_086_module_data_out[4] ,
    \sw_086_module_data_out[3] ,
    \sw_086_module_data_out[2] ,
    \sw_086_module_data_out[1] ,
    \sw_086_module_data_out[0] }));
 scanchain scanchain_087 (.clk_in(sw_086_clk_out),
    .clk_out(sw_087_clk_out),
    .data_in(sw_086_data_out),
    .data_out(sw_087_data_out),
    .latch_enable_in(sw_086_latch_out),
    .latch_enable_out(sw_087_latch_out),
    .scan_select_in(sw_086_scan_out),
    .scan_select_out(sw_087_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_087_module_data_in[7] ,
    \sw_087_module_data_in[6] ,
    \sw_087_module_data_in[5] ,
    \sw_087_module_data_in[4] ,
    \sw_087_module_data_in[3] ,
    \sw_087_module_data_in[2] ,
    \sw_087_module_data_in[1] ,
    \sw_087_module_data_in[0] }),
    .module_data_out({\sw_087_module_data_out[7] ,
    \sw_087_module_data_out[6] ,
    \sw_087_module_data_out[5] ,
    \sw_087_module_data_out[4] ,
    \sw_087_module_data_out[3] ,
    \sw_087_module_data_out[2] ,
    \sw_087_module_data_out[1] ,
    \sw_087_module_data_out[0] }));
 scanchain scanchain_088 (.clk_in(sw_087_clk_out),
    .clk_out(sw_088_clk_out),
    .data_in(sw_087_data_out),
    .data_out(sw_088_data_out),
    .latch_enable_in(sw_087_latch_out),
    .latch_enable_out(sw_088_latch_out),
    .scan_select_in(sw_087_scan_out),
    .scan_select_out(sw_088_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_088_module_data_in[7] ,
    \sw_088_module_data_in[6] ,
    \sw_088_module_data_in[5] ,
    \sw_088_module_data_in[4] ,
    \sw_088_module_data_in[3] ,
    \sw_088_module_data_in[2] ,
    \sw_088_module_data_in[1] ,
    \sw_088_module_data_in[0] }),
    .module_data_out({\sw_088_module_data_out[7] ,
    \sw_088_module_data_out[6] ,
    \sw_088_module_data_out[5] ,
    \sw_088_module_data_out[4] ,
    \sw_088_module_data_out[3] ,
    \sw_088_module_data_out[2] ,
    \sw_088_module_data_out[1] ,
    \sw_088_module_data_out[0] }));
 scanchain scanchain_089 (.clk_in(sw_088_clk_out),
    .clk_out(sw_089_clk_out),
    .data_in(sw_088_data_out),
    .data_out(sw_089_data_out),
    .latch_enable_in(sw_088_latch_out),
    .latch_enable_out(sw_089_latch_out),
    .scan_select_in(sw_088_scan_out),
    .scan_select_out(sw_089_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_089_module_data_in[7] ,
    \sw_089_module_data_in[6] ,
    \sw_089_module_data_in[5] ,
    \sw_089_module_data_in[4] ,
    \sw_089_module_data_in[3] ,
    \sw_089_module_data_in[2] ,
    \sw_089_module_data_in[1] ,
    \sw_089_module_data_in[0] }),
    .module_data_out({\sw_089_module_data_out[7] ,
    \sw_089_module_data_out[6] ,
    \sw_089_module_data_out[5] ,
    \sw_089_module_data_out[4] ,
    \sw_089_module_data_out[3] ,
    \sw_089_module_data_out[2] ,
    \sw_089_module_data_out[1] ,
    \sw_089_module_data_out[0] }));
 scanchain scanchain_090 (.clk_in(sw_089_clk_out),
    .clk_out(sw_090_clk_out),
    .data_in(sw_089_data_out),
    .data_out(sw_090_data_out),
    .latch_enable_in(sw_089_latch_out),
    .latch_enable_out(sw_090_latch_out),
    .scan_select_in(sw_089_scan_out),
    .scan_select_out(sw_090_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_090_module_data_in[7] ,
    \sw_090_module_data_in[6] ,
    \sw_090_module_data_in[5] ,
    \sw_090_module_data_in[4] ,
    \sw_090_module_data_in[3] ,
    \sw_090_module_data_in[2] ,
    \sw_090_module_data_in[1] ,
    \sw_090_module_data_in[0] }),
    .module_data_out({\sw_090_module_data_out[7] ,
    \sw_090_module_data_out[6] ,
    \sw_090_module_data_out[5] ,
    \sw_090_module_data_out[4] ,
    \sw_090_module_data_out[3] ,
    \sw_090_module_data_out[2] ,
    \sw_090_module_data_out[1] ,
    \sw_090_module_data_out[0] }));
 scanchain scanchain_091 (.clk_in(sw_090_clk_out),
    .clk_out(sw_091_clk_out),
    .data_in(sw_090_data_out),
    .data_out(sw_091_data_out),
    .latch_enable_in(sw_090_latch_out),
    .latch_enable_out(sw_091_latch_out),
    .scan_select_in(sw_090_scan_out),
    .scan_select_out(sw_091_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_091_module_data_in[7] ,
    \sw_091_module_data_in[6] ,
    \sw_091_module_data_in[5] ,
    \sw_091_module_data_in[4] ,
    \sw_091_module_data_in[3] ,
    \sw_091_module_data_in[2] ,
    \sw_091_module_data_in[1] ,
    \sw_091_module_data_in[0] }),
    .module_data_out({\sw_091_module_data_out[7] ,
    \sw_091_module_data_out[6] ,
    \sw_091_module_data_out[5] ,
    \sw_091_module_data_out[4] ,
    \sw_091_module_data_out[3] ,
    \sw_091_module_data_out[2] ,
    \sw_091_module_data_out[1] ,
    \sw_091_module_data_out[0] }));
 scanchain scanchain_092 (.clk_in(sw_091_clk_out),
    .clk_out(sw_092_clk_out),
    .data_in(sw_091_data_out),
    .data_out(sw_092_data_out),
    .latch_enable_in(sw_091_latch_out),
    .latch_enable_out(sw_092_latch_out),
    .scan_select_in(sw_091_scan_out),
    .scan_select_out(sw_092_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_092_module_data_in[7] ,
    \sw_092_module_data_in[6] ,
    \sw_092_module_data_in[5] ,
    \sw_092_module_data_in[4] ,
    \sw_092_module_data_in[3] ,
    \sw_092_module_data_in[2] ,
    \sw_092_module_data_in[1] ,
    \sw_092_module_data_in[0] }),
    .module_data_out({\sw_092_module_data_out[7] ,
    \sw_092_module_data_out[6] ,
    \sw_092_module_data_out[5] ,
    \sw_092_module_data_out[4] ,
    \sw_092_module_data_out[3] ,
    \sw_092_module_data_out[2] ,
    \sw_092_module_data_out[1] ,
    \sw_092_module_data_out[0] }));
 scanchain scanchain_093 (.clk_in(sw_092_clk_out),
    .clk_out(sw_093_clk_out),
    .data_in(sw_092_data_out),
    .data_out(sw_093_data_out),
    .latch_enable_in(sw_092_latch_out),
    .latch_enable_out(sw_093_latch_out),
    .scan_select_in(sw_092_scan_out),
    .scan_select_out(sw_093_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_093_module_data_in[7] ,
    \sw_093_module_data_in[6] ,
    \sw_093_module_data_in[5] ,
    \sw_093_module_data_in[4] ,
    \sw_093_module_data_in[3] ,
    \sw_093_module_data_in[2] ,
    \sw_093_module_data_in[1] ,
    \sw_093_module_data_in[0] }),
    .module_data_out({\sw_093_module_data_out[7] ,
    \sw_093_module_data_out[6] ,
    \sw_093_module_data_out[5] ,
    \sw_093_module_data_out[4] ,
    \sw_093_module_data_out[3] ,
    \sw_093_module_data_out[2] ,
    \sw_093_module_data_out[1] ,
    \sw_093_module_data_out[0] }));
 scanchain scanchain_094 (.clk_in(sw_093_clk_out),
    .clk_out(sw_094_clk_out),
    .data_in(sw_093_data_out),
    .data_out(sw_094_data_out),
    .latch_enable_in(sw_093_latch_out),
    .latch_enable_out(sw_094_latch_out),
    .scan_select_in(sw_093_scan_out),
    .scan_select_out(sw_094_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_094_module_data_in[7] ,
    \sw_094_module_data_in[6] ,
    \sw_094_module_data_in[5] ,
    \sw_094_module_data_in[4] ,
    \sw_094_module_data_in[3] ,
    \sw_094_module_data_in[2] ,
    \sw_094_module_data_in[1] ,
    \sw_094_module_data_in[0] }),
    .module_data_out({\sw_094_module_data_out[7] ,
    \sw_094_module_data_out[6] ,
    \sw_094_module_data_out[5] ,
    \sw_094_module_data_out[4] ,
    \sw_094_module_data_out[3] ,
    \sw_094_module_data_out[2] ,
    \sw_094_module_data_out[1] ,
    \sw_094_module_data_out[0] }));
 scanchain scanchain_095 (.clk_in(sw_094_clk_out),
    .clk_out(sw_095_clk_out),
    .data_in(sw_094_data_out),
    .data_out(sw_095_data_out),
    .latch_enable_in(sw_094_latch_out),
    .latch_enable_out(sw_095_latch_out),
    .scan_select_in(sw_094_scan_out),
    .scan_select_out(sw_095_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_095_module_data_in[7] ,
    \sw_095_module_data_in[6] ,
    \sw_095_module_data_in[5] ,
    \sw_095_module_data_in[4] ,
    \sw_095_module_data_in[3] ,
    \sw_095_module_data_in[2] ,
    \sw_095_module_data_in[1] ,
    \sw_095_module_data_in[0] }),
    .module_data_out({\sw_095_module_data_out[7] ,
    \sw_095_module_data_out[6] ,
    \sw_095_module_data_out[5] ,
    \sw_095_module_data_out[4] ,
    \sw_095_module_data_out[3] ,
    \sw_095_module_data_out[2] ,
    \sw_095_module_data_out[1] ,
    \sw_095_module_data_out[0] }));
 scanchain scanchain_096 (.clk_in(sw_095_clk_out),
    .clk_out(sw_096_clk_out),
    .data_in(sw_095_data_out),
    .data_out(sw_096_data_out),
    .latch_enable_in(sw_095_latch_out),
    .latch_enable_out(sw_096_latch_out),
    .scan_select_in(sw_095_scan_out),
    .scan_select_out(sw_096_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_096_module_data_in[7] ,
    \sw_096_module_data_in[6] ,
    \sw_096_module_data_in[5] ,
    \sw_096_module_data_in[4] ,
    \sw_096_module_data_in[3] ,
    \sw_096_module_data_in[2] ,
    \sw_096_module_data_in[1] ,
    \sw_096_module_data_in[0] }),
    .module_data_out({\sw_096_module_data_out[7] ,
    \sw_096_module_data_out[6] ,
    \sw_096_module_data_out[5] ,
    \sw_096_module_data_out[4] ,
    \sw_096_module_data_out[3] ,
    \sw_096_module_data_out[2] ,
    \sw_096_module_data_out[1] ,
    \sw_096_module_data_out[0] }));
 scanchain scanchain_097 (.clk_in(sw_096_clk_out),
    .clk_out(sw_097_clk_out),
    .data_in(sw_096_data_out),
    .data_out(sw_097_data_out),
    .latch_enable_in(sw_096_latch_out),
    .latch_enable_out(sw_097_latch_out),
    .scan_select_in(sw_096_scan_out),
    .scan_select_out(sw_097_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_097_module_data_in[7] ,
    \sw_097_module_data_in[6] ,
    \sw_097_module_data_in[5] ,
    \sw_097_module_data_in[4] ,
    \sw_097_module_data_in[3] ,
    \sw_097_module_data_in[2] ,
    \sw_097_module_data_in[1] ,
    \sw_097_module_data_in[0] }),
    .module_data_out({\sw_097_module_data_out[7] ,
    \sw_097_module_data_out[6] ,
    \sw_097_module_data_out[5] ,
    \sw_097_module_data_out[4] ,
    \sw_097_module_data_out[3] ,
    \sw_097_module_data_out[2] ,
    \sw_097_module_data_out[1] ,
    \sw_097_module_data_out[0] }));
 scanchain scanchain_098 (.clk_in(sw_097_clk_out),
    .clk_out(sw_098_clk_out),
    .data_in(sw_097_data_out),
    .data_out(sw_098_data_out),
    .latch_enable_in(sw_097_latch_out),
    .latch_enable_out(sw_098_latch_out),
    .scan_select_in(sw_097_scan_out),
    .scan_select_out(sw_098_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_098_module_data_in[7] ,
    \sw_098_module_data_in[6] ,
    \sw_098_module_data_in[5] ,
    \sw_098_module_data_in[4] ,
    \sw_098_module_data_in[3] ,
    \sw_098_module_data_in[2] ,
    \sw_098_module_data_in[1] ,
    \sw_098_module_data_in[0] }),
    .module_data_out({\sw_098_module_data_out[7] ,
    \sw_098_module_data_out[6] ,
    \sw_098_module_data_out[5] ,
    \sw_098_module_data_out[4] ,
    \sw_098_module_data_out[3] ,
    \sw_098_module_data_out[2] ,
    \sw_098_module_data_out[1] ,
    \sw_098_module_data_out[0] }));
 scanchain scanchain_099 (.clk_in(sw_098_clk_out),
    .clk_out(sw_099_clk_out),
    .data_in(sw_098_data_out),
    .data_out(sw_099_data_out),
    .latch_enable_in(sw_098_latch_out),
    .latch_enable_out(sw_099_latch_out),
    .scan_select_in(sw_098_scan_out),
    .scan_select_out(sw_099_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_099_module_data_in[7] ,
    \sw_099_module_data_in[6] ,
    \sw_099_module_data_in[5] ,
    \sw_099_module_data_in[4] ,
    \sw_099_module_data_in[3] ,
    \sw_099_module_data_in[2] ,
    \sw_099_module_data_in[1] ,
    \sw_099_module_data_in[0] }),
    .module_data_out({\sw_099_module_data_out[7] ,
    \sw_099_module_data_out[6] ,
    \sw_099_module_data_out[5] ,
    \sw_099_module_data_out[4] ,
    \sw_099_module_data_out[3] ,
    \sw_099_module_data_out[2] ,
    \sw_099_module_data_out[1] ,
    \sw_099_module_data_out[0] }));
 scanchain scanchain_100 (.clk_in(sw_099_clk_out),
    .clk_out(sw_100_clk_out),
    .data_in(sw_099_data_out),
    .data_out(sw_100_data_out),
    .latch_enable_in(sw_099_latch_out),
    .latch_enable_out(sw_100_latch_out),
    .scan_select_in(sw_099_scan_out),
    .scan_select_out(sw_100_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_100_module_data_in[7] ,
    \sw_100_module_data_in[6] ,
    \sw_100_module_data_in[5] ,
    \sw_100_module_data_in[4] ,
    \sw_100_module_data_in[3] ,
    \sw_100_module_data_in[2] ,
    \sw_100_module_data_in[1] ,
    \sw_100_module_data_in[0] }),
    .module_data_out({\sw_100_module_data_out[7] ,
    \sw_100_module_data_out[6] ,
    \sw_100_module_data_out[5] ,
    \sw_100_module_data_out[4] ,
    \sw_100_module_data_out[3] ,
    \sw_100_module_data_out[2] ,
    \sw_100_module_data_out[1] ,
    \sw_100_module_data_out[0] }));
 scanchain scanchain_101 (.clk_in(sw_100_clk_out),
    .clk_out(sw_101_clk_out),
    .data_in(sw_100_data_out),
    .data_out(sw_101_data_out),
    .latch_enable_in(sw_100_latch_out),
    .latch_enable_out(sw_101_latch_out),
    .scan_select_in(sw_100_scan_out),
    .scan_select_out(sw_101_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_101_module_data_in[7] ,
    \sw_101_module_data_in[6] ,
    \sw_101_module_data_in[5] ,
    \sw_101_module_data_in[4] ,
    \sw_101_module_data_in[3] ,
    \sw_101_module_data_in[2] ,
    \sw_101_module_data_in[1] ,
    \sw_101_module_data_in[0] }),
    .module_data_out({\sw_101_module_data_out[7] ,
    \sw_101_module_data_out[6] ,
    \sw_101_module_data_out[5] ,
    \sw_101_module_data_out[4] ,
    \sw_101_module_data_out[3] ,
    \sw_101_module_data_out[2] ,
    \sw_101_module_data_out[1] ,
    \sw_101_module_data_out[0] }));
 scanchain scanchain_102 (.clk_in(sw_101_clk_out),
    .clk_out(sw_102_clk_out),
    .data_in(sw_101_data_out),
    .data_out(sw_102_data_out),
    .latch_enable_in(sw_101_latch_out),
    .latch_enable_out(sw_102_latch_out),
    .scan_select_in(sw_101_scan_out),
    .scan_select_out(sw_102_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_102_module_data_in[7] ,
    \sw_102_module_data_in[6] ,
    \sw_102_module_data_in[5] ,
    \sw_102_module_data_in[4] ,
    \sw_102_module_data_in[3] ,
    \sw_102_module_data_in[2] ,
    \sw_102_module_data_in[1] ,
    \sw_102_module_data_in[0] }),
    .module_data_out({\sw_102_module_data_out[7] ,
    \sw_102_module_data_out[6] ,
    \sw_102_module_data_out[5] ,
    \sw_102_module_data_out[4] ,
    \sw_102_module_data_out[3] ,
    \sw_102_module_data_out[2] ,
    \sw_102_module_data_out[1] ,
    \sw_102_module_data_out[0] }));
 scanchain scanchain_103 (.clk_in(sw_102_clk_out),
    .clk_out(sw_103_clk_out),
    .data_in(sw_102_data_out),
    .data_out(sw_103_data_out),
    .latch_enable_in(sw_102_latch_out),
    .latch_enable_out(sw_103_latch_out),
    .scan_select_in(sw_102_scan_out),
    .scan_select_out(sw_103_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_103_module_data_in[7] ,
    \sw_103_module_data_in[6] ,
    \sw_103_module_data_in[5] ,
    \sw_103_module_data_in[4] ,
    \sw_103_module_data_in[3] ,
    \sw_103_module_data_in[2] ,
    \sw_103_module_data_in[1] ,
    \sw_103_module_data_in[0] }),
    .module_data_out({\sw_103_module_data_out[7] ,
    \sw_103_module_data_out[6] ,
    \sw_103_module_data_out[5] ,
    \sw_103_module_data_out[4] ,
    \sw_103_module_data_out[3] ,
    \sw_103_module_data_out[2] ,
    \sw_103_module_data_out[1] ,
    \sw_103_module_data_out[0] }));
 scanchain scanchain_104 (.clk_in(sw_103_clk_out),
    .clk_out(sw_104_clk_out),
    .data_in(sw_103_data_out),
    .data_out(sw_104_data_out),
    .latch_enable_in(sw_103_latch_out),
    .latch_enable_out(sw_104_latch_out),
    .scan_select_in(sw_103_scan_out),
    .scan_select_out(sw_104_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_104_module_data_in[7] ,
    \sw_104_module_data_in[6] ,
    \sw_104_module_data_in[5] ,
    \sw_104_module_data_in[4] ,
    \sw_104_module_data_in[3] ,
    \sw_104_module_data_in[2] ,
    \sw_104_module_data_in[1] ,
    \sw_104_module_data_in[0] }),
    .module_data_out({\sw_104_module_data_out[7] ,
    \sw_104_module_data_out[6] ,
    \sw_104_module_data_out[5] ,
    \sw_104_module_data_out[4] ,
    \sw_104_module_data_out[3] ,
    \sw_104_module_data_out[2] ,
    \sw_104_module_data_out[1] ,
    \sw_104_module_data_out[0] }));
 scanchain scanchain_105 (.clk_in(sw_104_clk_out),
    .clk_out(sw_105_clk_out),
    .data_in(sw_104_data_out),
    .data_out(sw_105_data_out),
    .latch_enable_in(sw_104_latch_out),
    .latch_enable_out(sw_105_latch_out),
    .scan_select_in(sw_104_scan_out),
    .scan_select_out(sw_105_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_105_module_data_in[7] ,
    \sw_105_module_data_in[6] ,
    \sw_105_module_data_in[5] ,
    \sw_105_module_data_in[4] ,
    \sw_105_module_data_in[3] ,
    \sw_105_module_data_in[2] ,
    \sw_105_module_data_in[1] ,
    \sw_105_module_data_in[0] }),
    .module_data_out({\sw_105_module_data_out[7] ,
    \sw_105_module_data_out[6] ,
    \sw_105_module_data_out[5] ,
    \sw_105_module_data_out[4] ,
    \sw_105_module_data_out[3] ,
    \sw_105_module_data_out[2] ,
    \sw_105_module_data_out[1] ,
    \sw_105_module_data_out[0] }));
 scanchain scanchain_106 (.clk_in(sw_105_clk_out),
    .clk_out(sw_106_clk_out),
    .data_in(sw_105_data_out),
    .data_out(sw_106_data_out),
    .latch_enable_in(sw_105_latch_out),
    .latch_enable_out(sw_106_latch_out),
    .scan_select_in(sw_105_scan_out),
    .scan_select_out(sw_106_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_106_module_data_in[7] ,
    \sw_106_module_data_in[6] ,
    \sw_106_module_data_in[5] ,
    \sw_106_module_data_in[4] ,
    \sw_106_module_data_in[3] ,
    \sw_106_module_data_in[2] ,
    \sw_106_module_data_in[1] ,
    \sw_106_module_data_in[0] }),
    .module_data_out({\sw_106_module_data_out[7] ,
    \sw_106_module_data_out[6] ,
    \sw_106_module_data_out[5] ,
    \sw_106_module_data_out[4] ,
    \sw_106_module_data_out[3] ,
    \sw_106_module_data_out[2] ,
    \sw_106_module_data_out[1] ,
    \sw_106_module_data_out[0] }));
 scanchain scanchain_107 (.clk_in(sw_106_clk_out),
    .clk_out(sw_107_clk_out),
    .data_in(sw_106_data_out),
    .data_out(sw_107_data_out),
    .latch_enable_in(sw_106_latch_out),
    .latch_enable_out(sw_107_latch_out),
    .scan_select_in(sw_106_scan_out),
    .scan_select_out(sw_107_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_107_module_data_in[7] ,
    \sw_107_module_data_in[6] ,
    \sw_107_module_data_in[5] ,
    \sw_107_module_data_in[4] ,
    \sw_107_module_data_in[3] ,
    \sw_107_module_data_in[2] ,
    \sw_107_module_data_in[1] ,
    \sw_107_module_data_in[0] }),
    .module_data_out({\sw_107_module_data_out[7] ,
    \sw_107_module_data_out[6] ,
    \sw_107_module_data_out[5] ,
    \sw_107_module_data_out[4] ,
    \sw_107_module_data_out[3] ,
    \sw_107_module_data_out[2] ,
    \sw_107_module_data_out[1] ,
    \sw_107_module_data_out[0] }));
 scanchain scanchain_108 (.clk_in(sw_107_clk_out),
    .clk_out(sw_108_clk_out),
    .data_in(sw_107_data_out),
    .data_out(sw_108_data_out),
    .latch_enable_in(sw_107_latch_out),
    .latch_enable_out(sw_108_latch_out),
    .scan_select_in(sw_107_scan_out),
    .scan_select_out(sw_108_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_108_module_data_in[7] ,
    \sw_108_module_data_in[6] ,
    \sw_108_module_data_in[5] ,
    \sw_108_module_data_in[4] ,
    \sw_108_module_data_in[3] ,
    \sw_108_module_data_in[2] ,
    \sw_108_module_data_in[1] ,
    \sw_108_module_data_in[0] }),
    .module_data_out({\sw_108_module_data_out[7] ,
    \sw_108_module_data_out[6] ,
    \sw_108_module_data_out[5] ,
    \sw_108_module_data_out[4] ,
    \sw_108_module_data_out[3] ,
    \sw_108_module_data_out[2] ,
    \sw_108_module_data_out[1] ,
    \sw_108_module_data_out[0] }));
 scanchain scanchain_109 (.clk_in(sw_108_clk_out),
    .clk_out(sw_109_clk_out),
    .data_in(sw_108_data_out),
    .data_out(sw_109_data_out),
    .latch_enable_in(sw_108_latch_out),
    .latch_enable_out(sw_109_latch_out),
    .scan_select_in(sw_108_scan_out),
    .scan_select_out(sw_109_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_109_module_data_in[7] ,
    \sw_109_module_data_in[6] ,
    \sw_109_module_data_in[5] ,
    \sw_109_module_data_in[4] ,
    \sw_109_module_data_in[3] ,
    \sw_109_module_data_in[2] ,
    \sw_109_module_data_in[1] ,
    \sw_109_module_data_in[0] }),
    .module_data_out({\sw_109_module_data_out[7] ,
    \sw_109_module_data_out[6] ,
    \sw_109_module_data_out[5] ,
    \sw_109_module_data_out[4] ,
    \sw_109_module_data_out[3] ,
    \sw_109_module_data_out[2] ,
    \sw_109_module_data_out[1] ,
    \sw_109_module_data_out[0] }));
 scanchain scanchain_110 (.clk_in(sw_109_clk_out),
    .clk_out(sw_110_clk_out),
    .data_in(sw_109_data_out),
    .data_out(sw_110_data_out),
    .latch_enable_in(sw_109_latch_out),
    .latch_enable_out(sw_110_latch_out),
    .scan_select_in(sw_109_scan_out),
    .scan_select_out(sw_110_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_110_module_data_in[7] ,
    \sw_110_module_data_in[6] ,
    \sw_110_module_data_in[5] ,
    \sw_110_module_data_in[4] ,
    \sw_110_module_data_in[3] ,
    \sw_110_module_data_in[2] ,
    \sw_110_module_data_in[1] ,
    \sw_110_module_data_in[0] }),
    .module_data_out({\sw_110_module_data_out[7] ,
    \sw_110_module_data_out[6] ,
    \sw_110_module_data_out[5] ,
    \sw_110_module_data_out[4] ,
    \sw_110_module_data_out[3] ,
    \sw_110_module_data_out[2] ,
    \sw_110_module_data_out[1] ,
    \sw_110_module_data_out[0] }));
 scanchain scanchain_111 (.clk_in(sw_110_clk_out),
    .clk_out(sw_111_clk_out),
    .data_in(sw_110_data_out),
    .data_out(sw_111_data_out),
    .latch_enable_in(sw_110_latch_out),
    .latch_enable_out(sw_111_latch_out),
    .scan_select_in(sw_110_scan_out),
    .scan_select_out(sw_111_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_111_module_data_in[7] ,
    \sw_111_module_data_in[6] ,
    \sw_111_module_data_in[5] ,
    \sw_111_module_data_in[4] ,
    \sw_111_module_data_in[3] ,
    \sw_111_module_data_in[2] ,
    \sw_111_module_data_in[1] ,
    \sw_111_module_data_in[0] }),
    .module_data_out({\sw_111_module_data_out[7] ,
    \sw_111_module_data_out[6] ,
    \sw_111_module_data_out[5] ,
    \sw_111_module_data_out[4] ,
    \sw_111_module_data_out[3] ,
    \sw_111_module_data_out[2] ,
    \sw_111_module_data_out[1] ,
    \sw_111_module_data_out[0] }));
 scanchain scanchain_112 (.clk_in(sw_111_clk_out),
    .clk_out(sw_112_clk_out),
    .data_in(sw_111_data_out),
    .data_out(sw_112_data_out),
    .latch_enable_in(sw_111_latch_out),
    .latch_enable_out(sw_112_latch_out),
    .scan_select_in(sw_111_scan_out),
    .scan_select_out(sw_112_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_112_module_data_in[7] ,
    \sw_112_module_data_in[6] ,
    \sw_112_module_data_in[5] ,
    \sw_112_module_data_in[4] ,
    \sw_112_module_data_in[3] ,
    \sw_112_module_data_in[2] ,
    \sw_112_module_data_in[1] ,
    \sw_112_module_data_in[0] }),
    .module_data_out({\sw_112_module_data_out[7] ,
    \sw_112_module_data_out[6] ,
    \sw_112_module_data_out[5] ,
    \sw_112_module_data_out[4] ,
    \sw_112_module_data_out[3] ,
    \sw_112_module_data_out[2] ,
    \sw_112_module_data_out[1] ,
    \sw_112_module_data_out[0] }));
 scanchain scanchain_113 (.clk_in(sw_112_clk_out),
    .clk_out(sw_113_clk_out),
    .data_in(sw_112_data_out),
    .data_out(sw_113_data_out),
    .latch_enable_in(sw_112_latch_out),
    .latch_enable_out(sw_113_latch_out),
    .scan_select_in(sw_112_scan_out),
    .scan_select_out(sw_113_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_113_module_data_in[7] ,
    \sw_113_module_data_in[6] ,
    \sw_113_module_data_in[5] ,
    \sw_113_module_data_in[4] ,
    \sw_113_module_data_in[3] ,
    \sw_113_module_data_in[2] ,
    \sw_113_module_data_in[1] ,
    \sw_113_module_data_in[0] }),
    .module_data_out({\sw_113_module_data_out[7] ,
    \sw_113_module_data_out[6] ,
    \sw_113_module_data_out[5] ,
    \sw_113_module_data_out[4] ,
    \sw_113_module_data_out[3] ,
    \sw_113_module_data_out[2] ,
    \sw_113_module_data_out[1] ,
    \sw_113_module_data_out[0] }));
 scanchain scanchain_114 (.clk_in(sw_113_clk_out),
    .clk_out(sw_114_clk_out),
    .data_in(sw_113_data_out),
    .data_out(sw_114_data_out),
    .latch_enable_in(sw_113_latch_out),
    .latch_enable_out(sw_114_latch_out),
    .scan_select_in(sw_113_scan_out),
    .scan_select_out(sw_114_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_114_module_data_in[7] ,
    \sw_114_module_data_in[6] ,
    \sw_114_module_data_in[5] ,
    \sw_114_module_data_in[4] ,
    \sw_114_module_data_in[3] ,
    \sw_114_module_data_in[2] ,
    \sw_114_module_data_in[1] ,
    \sw_114_module_data_in[0] }),
    .module_data_out({\sw_114_module_data_out[7] ,
    \sw_114_module_data_out[6] ,
    \sw_114_module_data_out[5] ,
    \sw_114_module_data_out[4] ,
    \sw_114_module_data_out[3] ,
    \sw_114_module_data_out[2] ,
    \sw_114_module_data_out[1] ,
    \sw_114_module_data_out[0] }));
 scanchain scanchain_115 (.clk_in(sw_114_clk_out),
    .clk_out(sw_115_clk_out),
    .data_in(sw_114_data_out),
    .data_out(sw_115_data_out),
    .latch_enable_in(sw_114_latch_out),
    .latch_enable_out(sw_115_latch_out),
    .scan_select_in(sw_114_scan_out),
    .scan_select_out(sw_115_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_115_module_data_in[7] ,
    \sw_115_module_data_in[6] ,
    \sw_115_module_data_in[5] ,
    \sw_115_module_data_in[4] ,
    \sw_115_module_data_in[3] ,
    \sw_115_module_data_in[2] ,
    \sw_115_module_data_in[1] ,
    \sw_115_module_data_in[0] }),
    .module_data_out({\sw_115_module_data_out[7] ,
    \sw_115_module_data_out[6] ,
    \sw_115_module_data_out[5] ,
    \sw_115_module_data_out[4] ,
    \sw_115_module_data_out[3] ,
    \sw_115_module_data_out[2] ,
    \sw_115_module_data_out[1] ,
    \sw_115_module_data_out[0] }));
 scanchain scanchain_116 (.clk_in(sw_115_clk_out),
    .clk_out(sw_116_clk_out),
    .data_in(sw_115_data_out),
    .data_out(sw_116_data_out),
    .latch_enable_in(sw_115_latch_out),
    .latch_enable_out(sw_116_latch_out),
    .scan_select_in(sw_115_scan_out),
    .scan_select_out(sw_116_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_116_module_data_in[7] ,
    \sw_116_module_data_in[6] ,
    \sw_116_module_data_in[5] ,
    \sw_116_module_data_in[4] ,
    \sw_116_module_data_in[3] ,
    \sw_116_module_data_in[2] ,
    \sw_116_module_data_in[1] ,
    \sw_116_module_data_in[0] }),
    .module_data_out({\sw_116_module_data_out[7] ,
    \sw_116_module_data_out[6] ,
    \sw_116_module_data_out[5] ,
    \sw_116_module_data_out[4] ,
    \sw_116_module_data_out[3] ,
    \sw_116_module_data_out[2] ,
    \sw_116_module_data_out[1] ,
    \sw_116_module_data_out[0] }));
 scanchain scanchain_117 (.clk_in(sw_116_clk_out),
    .clk_out(sw_117_clk_out),
    .data_in(sw_116_data_out),
    .data_out(sw_117_data_out),
    .latch_enable_in(sw_116_latch_out),
    .latch_enable_out(sw_117_latch_out),
    .scan_select_in(sw_116_scan_out),
    .scan_select_out(sw_117_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_117_module_data_in[7] ,
    \sw_117_module_data_in[6] ,
    \sw_117_module_data_in[5] ,
    \sw_117_module_data_in[4] ,
    \sw_117_module_data_in[3] ,
    \sw_117_module_data_in[2] ,
    \sw_117_module_data_in[1] ,
    \sw_117_module_data_in[0] }),
    .module_data_out({\sw_117_module_data_out[7] ,
    \sw_117_module_data_out[6] ,
    \sw_117_module_data_out[5] ,
    \sw_117_module_data_out[4] ,
    \sw_117_module_data_out[3] ,
    \sw_117_module_data_out[2] ,
    \sw_117_module_data_out[1] ,
    \sw_117_module_data_out[0] }));
 scanchain scanchain_118 (.clk_in(sw_117_clk_out),
    .clk_out(sw_118_clk_out),
    .data_in(sw_117_data_out),
    .data_out(sw_118_data_out),
    .latch_enable_in(sw_117_latch_out),
    .latch_enable_out(sw_118_latch_out),
    .scan_select_in(sw_117_scan_out),
    .scan_select_out(sw_118_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_118_module_data_in[7] ,
    \sw_118_module_data_in[6] ,
    \sw_118_module_data_in[5] ,
    \sw_118_module_data_in[4] ,
    \sw_118_module_data_in[3] ,
    \sw_118_module_data_in[2] ,
    \sw_118_module_data_in[1] ,
    \sw_118_module_data_in[0] }),
    .module_data_out({\sw_118_module_data_out[7] ,
    \sw_118_module_data_out[6] ,
    \sw_118_module_data_out[5] ,
    \sw_118_module_data_out[4] ,
    \sw_118_module_data_out[3] ,
    \sw_118_module_data_out[2] ,
    \sw_118_module_data_out[1] ,
    \sw_118_module_data_out[0] }));
 scanchain scanchain_119 (.clk_in(sw_118_clk_out),
    .clk_out(sw_119_clk_out),
    .data_in(sw_118_data_out),
    .data_out(sw_119_data_out),
    .latch_enable_in(sw_118_latch_out),
    .latch_enable_out(sw_119_latch_out),
    .scan_select_in(sw_118_scan_out),
    .scan_select_out(sw_119_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_119_module_data_in[7] ,
    \sw_119_module_data_in[6] ,
    \sw_119_module_data_in[5] ,
    \sw_119_module_data_in[4] ,
    \sw_119_module_data_in[3] ,
    \sw_119_module_data_in[2] ,
    \sw_119_module_data_in[1] ,
    \sw_119_module_data_in[0] }),
    .module_data_out({\sw_119_module_data_out[7] ,
    \sw_119_module_data_out[6] ,
    \sw_119_module_data_out[5] ,
    \sw_119_module_data_out[4] ,
    \sw_119_module_data_out[3] ,
    \sw_119_module_data_out[2] ,
    \sw_119_module_data_out[1] ,
    \sw_119_module_data_out[0] }));
 scanchain scanchain_120 (.clk_in(sw_119_clk_out),
    .clk_out(sw_120_clk_out),
    .data_in(sw_119_data_out),
    .data_out(sw_120_data_out),
    .latch_enable_in(sw_119_latch_out),
    .latch_enable_out(sw_120_latch_out),
    .scan_select_in(sw_119_scan_out),
    .scan_select_out(sw_120_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_120_module_data_in[7] ,
    \sw_120_module_data_in[6] ,
    \sw_120_module_data_in[5] ,
    \sw_120_module_data_in[4] ,
    \sw_120_module_data_in[3] ,
    \sw_120_module_data_in[2] ,
    \sw_120_module_data_in[1] ,
    \sw_120_module_data_in[0] }),
    .module_data_out({\sw_120_module_data_out[7] ,
    \sw_120_module_data_out[6] ,
    \sw_120_module_data_out[5] ,
    \sw_120_module_data_out[4] ,
    \sw_120_module_data_out[3] ,
    \sw_120_module_data_out[2] ,
    \sw_120_module_data_out[1] ,
    \sw_120_module_data_out[0] }));
 scanchain scanchain_121 (.clk_in(sw_120_clk_out),
    .clk_out(sw_121_clk_out),
    .data_in(sw_120_data_out),
    .data_out(sw_121_data_out),
    .latch_enable_in(sw_120_latch_out),
    .latch_enable_out(sw_121_latch_out),
    .scan_select_in(sw_120_scan_out),
    .scan_select_out(sw_121_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_121_module_data_in[7] ,
    \sw_121_module_data_in[6] ,
    \sw_121_module_data_in[5] ,
    \sw_121_module_data_in[4] ,
    \sw_121_module_data_in[3] ,
    \sw_121_module_data_in[2] ,
    \sw_121_module_data_in[1] ,
    \sw_121_module_data_in[0] }),
    .module_data_out({\sw_121_module_data_out[7] ,
    \sw_121_module_data_out[6] ,
    \sw_121_module_data_out[5] ,
    \sw_121_module_data_out[4] ,
    \sw_121_module_data_out[3] ,
    \sw_121_module_data_out[2] ,
    \sw_121_module_data_out[1] ,
    \sw_121_module_data_out[0] }));
 scanchain scanchain_122 (.clk_in(sw_121_clk_out),
    .clk_out(sw_122_clk_out),
    .data_in(sw_121_data_out),
    .data_out(sw_122_data_out),
    .latch_enable_in(sw_121_latch_out),
    .latch_enable_out(sw_122_latch_out),
    .scan_select_in(sw_121_scan_out),
    .scan_select_out(sw_122_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_122_module_data_in[7] ,
    \sw_122_module_data_in[6] ,
    \sw_122_module_data_in[5] ,
    \sw_122_module_data_in[4] ,
    \sw_122_module_data_in[3] ,
    \sw_122_module_data_in[2] ,
    \sw_122_module_data_in[1] ,
    \sw_122_module_data_in[0] }),
    .module_data_out({\sw_122_module_data_out[7] ,
    \sw_122_module_data_out[6] ,
    \sw_122_module_data_out[5] ,
    \sw_122_module_data_out[4] ,
    \sw_122_module_data_out[3] ,
    \sw_122_module_data_out[2] ,
    \sw_122_module_data_out[1] ,
    \sw_122_module_data_out[0] }));
 scanchain scanchain_123 (.clk_in(sw_122_clk_out),
    .clk_out(sw_123_clk_out),
    .data_in(sw_122_data_out),
    .data_out(sw_123_data_out),
    .latch_enable_in(sw_122_latch_out),
    .latch_enable_out(sw_123_latch_out),
    .scan_select_in(sw_122_scan_out),
    .scan_select_out(sw_123_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_123_module_data_in[7] ,
    \sw_123_module_data_in[6] ,
    \sw_123_module_data_in[5] ,
    \sw_123_module_data_in[4] ,
    \sw_123_module_data_in[3] ,
    \sw_123_module_data_in[2] ,
    \sw_123_module_data_in[1] ,
    \sw_123_module_data_in[0] }),
    .module_data_out({\sw_123_module_data_out[7] ,
    \sw_123_module_data_out[6] ,
    \sw_123_module_data_out[5] ,
    \sw_123_module_data_out[4] ,
    \sw_123_module_data_out[3] ,
    \sw_123_module_data_out[2] ,
    \sw_123_module_data_out[1] ,
    \sw_123_module_data_out[0] }));
 scanchain scanchain_124 (.clk_in(sw_123_clk_out),
    .clk_out(sw_124_clk_out),
    .data_in(sw_123_data_out),
    .data_out(sw_124_data_out),
    .latch_enable_in(sw_123_latch_out),
    .latch_enable_out(sw_124_latch_out),
    .scan_select_in(sw_123_scan_out),
    .scan_select_out(sw_124_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_124_module_data_in[7] ,
    \sw_124_module_data_in[6] ,
    \sw_124_module_data_in[5] ,
    \sw_124_module_data_in[4] ,
    \sw_124_module_data_in[3] ,
    \sw_124_module_data_in[2] ,
    \sw_124_module_data_in[1] ,
    \sw_124_module_data_in[0] }),
    .module_data_out({\sw_124_module_data_out[7] ,
    \sw_124_module_data_out[6] ,
    \sw_124_module_data_out[5] ,
    \sw_124_module_data_out[4] ,
    \sw_124_module_data_out[3] ,
    \sw_124_module_data_out[2] ,
    \sw_124_module_data_out[1] ,
    \sw_124_module_data_out[0] }));
 scanchain scanchain_125 (.clk_in(sw_124_clk_out),
    .clk_out(sw_125_clk_out),
    .data_in(sw_124_data_out),
    .data_out(sw_125_data_out),
    .latch_enable_in(sw_124_latch_out),
    .latch_enable_out(sw_125_latch_out),
    .scan_select_in(sw_124_scan_out),
    .scan_select_out(sw_125_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_125_module_data_in[7] ,
    \sw_125_module_data_in[6] ,
    \sw_125_module_data_in[5] ,
    \sw_125_module_data_in[4] ,
    \sw_125_module_data_in[3] ,
    \sw_125_module_data_in[2] ,
    \sw_125_module_data_in[1] ,
    \sw_125_module_data_in[0] }),
    .module_data_out({\sw_125_module_data_out[7] ,
    \sw_125_module_data_out[6] ,
    \sw_125_module_data_out[5] ,
    \sw_125_module_data_out[4] ,
    \sw_125_module_data_out[3] ,
    \sw_125_module_data_out[2] ,
    \sw_125_module_data_out[1] ,
    \sw_125_module_data_out[0] }));
 scanchain scanchain_126 (.clk_in(sw_125_clk_out),
    .clk_out(sw_126_clk_out),
    .data_in(sw_125_data_out),
    .data_out(sw_126_data_out),
    .latch_enable_in(sw_125_latch_out),
    .latch_enable_out(sw_126_latch_out),
    .scan_select_in(sw_125_scan_out),
    .scan_select_out(sw_126_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_126_module_data_in[7] ,
    \sw_126_module_data_in[6] ,
    \sw_126_module_data_in[5] ,
    \sw_126_module_data_in[4] ,
    \sw_126_module_data_in[3] ,
    \sw_126_module_data_in[2] ,
    \sw_126_module_data_in[1] ,
    \sw_126_module_data_in[0] }),
    .module_data_out({\sw_126_module_data_out[7] ,
    \sw_126_module_data_out[6] ,
    \sw_126_module_data_out[5] ,
    \sw_126_module_data_out[4] ,
    \sw_126_module_data_out[3] ,
    \sw_126_module_data_out[2] ,
    \sw_126_module_data_out[1] ,
    \sw_126_module_data_out[0] }));
 scanchain scanchain_127 (.clk_in(sw_126_clk_out),
    .clk_out(sw_127_clk_out),
    .data_in(sw_126_data_out),
    .data_out(sw_127_data_out),
    .latch_enable_in(sw_126_latch_out),
    .latch_enable_out(sw_127_latch_out),
    .scan_select_in(sw_126_scan_out),
    .scan_select_out(sw_127_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_127_module_data_in[7] ,
    \sw_127_module_data_in[6] ,
    \sw_127_module_data_in[5] ,
    \sw_127_module_data_in[4] ,
    \sw_127_module_data_in[3] ,
    \sw_127_module_data_in[2] ,
    \sw_127_module_data_in[1] ,
    \sw_127_module_data_in[0] }),
    .module_data_out({\sw_127_module_data_out[7] ,
    \sw_127_module_data_out[6] ,
    \sw_127_module_data_out[5] ,
    \sw_127_module_data_out[4] ,
    \sw_127_module_data_out[3] ,
    \sw_127_module_data_out[2] ,
    \sw_127_module_data_out[1] ,
    \sw_127_module_data_out[0] }));
 scanchain scanchain_128 (.clk_in(sw_127_clk_out),
    .clk_out(sw_128_clk_out),
    .data_in(sw_127_data_out),
    .data_out(sw_128_data_out),
    .latch_enable_in(sw_127_latch_out),
    .latch_enable_out(sw_128_latch_out),
    .scan_select_in(sw_127_scan_out),
    .scan_select_out(sw_128_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_128_module_data_in[7] ,
    \sw_128_module_data_in[6] ,
    \sw_128_module_data_in[5] ,
    \sw_128_module_data_in[4] ,
    \sw_128_module_data_in[3] ,
    \sw_128_module_data_in[2] ,
    \sw_128_module_data_in[1] ,
    \sw_128_module_data_in[0] }),
    .module_data_out({\sw_128_module_data_out[7] ,
    \sw_128_module_data_out[6] ,
    \sw_128_module_data_out[5] ,
    \sw_128_module_data_out[4] ,
    \sw_128_module_data_out[3] ,
    \sw_128_module_data_out[2] ,
    \sw_128_module_data_out[1] ,
    \sw_128_module_data_out[0] }));
 scanchain scanchain_129 (.clk_in(sw_128_clk_out),
    .clk_out(sw_129_clk_out),
    .data_in(sw_128_data_out),
    .data_out(sw_129_data_out),
    .latch_enable_in(sw_128_latch_out),
    .latch_enable_out(sw_129_latch_out),
    .scan_select_in(sw_128_scan_out),
    .scan_select_out(sw_129_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_129_module_data_in[7] ,
    \sw_129_module_data_in[6] ,
    \sw_129_module_data_in[5] ,
    \sw_129_module_data_in[4] ,
    \sw_129_module_data_in[3] ,
    \sw_129_module_data_in[2] ,
    \sw_129_module_data_in[1] ,
    \sw_129_module_data_in[0] }),
    .module_data_out({\sw_129_module_data_out[7] ,
    \sw_129_module_data_out[6] ,
    \sw_129_module_data_out[5] ,
    \sw_129_module_data_out[4] ,
    \sw_129_module_data_out[3] ,
    \sw_129_module_data_out[2] ,
    \sw_129_module_data_out[1] ,
    \sw_129_module_data_out[0] }));
 scanchain scanchain_130 (.clk_in(sw_129_clk_out),
    .clk_out(sw_130_clk_out),
    .data_in(sw_129_data_out),
    .data_out(sw_130_data_out),
    .latch_enable_in(sw_129_latch_out),
    .latch_enable_out(sw_130_latch_out),
    .scan_select_in(sw_129_scan_out),
    .scan_select_out(sw_130_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_130_module_data_in[7] ,
    \sw_130_module_data_in[6] ,
    \sw_130_module_data_in[5] ,
    \sw_130_module_data_in[4] ,
    \sw_130_module_data_in[3] ,
    \sw_130_module_data_in[2] ,
    \sw_130_module_data_in[1] ,
    \sw_130_module_data_in[0] }),
    .module_data_out({\sw_130_module_data_out[7] ,
    \sw_130_module_data_out[6] ,
    \sw_130_module_data_out[5] ,
    \sw_130_module_data_out[4] ,
    \sw_130_module_data_out[3] ,
    \sw_130_module_data_out[2] ,
    \sw_130_module_data_out[1] ,
    \sw_130_module_data_out[0] }));
 scanchain scanchain_131 (.clk_in(sw_130_clk_out),
    .clk_out(sw_131_clk_out),
    .data_in(sw_130_data_out),
    .data_out(sw_131_data_out),
    .latch_enable_in(sw_130_latch_out),
    .latch_enable_out(sw_131_latch_out),
    .scan_select_in(sw_130_scan_out),
    .scan_select_out(sw_131_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_131_module_data_in[7] ,
    \sw_131_module_data_in[6] ,
    \sw_131_module_data_in[5] ,
    \sw_131_module_data_in[4] ,
    \sw_131_module_data_in[3] ,
    \sw_131_module_data_in[2] ,
    \sw_131_module_data_in[1] ,
    \sw_131_module_data_in[0] }),
    .module_data_out({\sw_131_module_data_out[7] ,
    \sw_131_module_data_out[6] ,
    \sw_131_module_data_out[5] ,
    \sw_131_module_data_out[4] ,
    \sw_131_module_data_out[3] ,
    \sw_131_module_data_out[2] ,
    \sw_131_module_data_out[1] ,
    \sw_131_module_data_out[0] }));
 scanchain scanchain_132 (.clk_in(sw_131_clk_out),
    .clk_out(sw_132_clk_out),
    .data_in(sw_131_data_out),
    .data_out(sw_132_data_out),
    .latch_enable_in(sw_131_latch_out),
    .latch_enable_out(sw_132_latch_out),
    .scan_select_in(sw_131_scan_out),
    .scan_select_out(sw_132_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_132_module_data_in[7] ,
    \sw_132_module_data_in[6] ,
    \sw_132_module_data_in[5] ,
    \sw_132_module_data_in[4] ,
    \sw_132_module_data_in[3] ,
    \sw_132_module_data_in[2] ,
    \sw_132_module_data_in[1] ,
    \sw_132_module_data_in[0] }),
    .module_data_out({\sw_132_module_data_out[7] ,
    \sw_132_module_data_out[6] ,
    \sw_132_module_data_out[5] ,
    \sw_132_module_data_out[4] ,
    \sw_132_module_data_out[3] ,
    \sw_132_module_data_out[2] ,
    \sw_132_module_data_out[1] ,
    \sw_132_module_data_out[0] }));
 scanchain scanchain_133 (.clk_in(sw_132_clk_out),
    .clk_out(sw_133_clk_out),
    .data_in(sw_132_data_out),
    .data_out(sw_133_data_out),
    .latch_enable_in(sw_132_latch_out),
    .latch_enable_out(sw_133_latch_out),
    .scan_select_in(sw_132_scan_out),
    .scan_select_out(sw_133_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_133_module_data_in[7] ,
    \sw_133_module_data_in[6] ,
    \sw_133_module_data_in[5] ,
    \sw_133_module_data_in[4] ,
    \sw_133_module_data_in[3] ,
    \sw_133_module_data_in[2] ,
    \sw_133_module_data_in[1] ,
    \sw_133_module_data_in[0] }),
    .module_data_out({\sw_133_module_data_out[7] ,
    \sw_133_module_data_out[6] ,
    \sw_133_module_data_out[5] ,
    \sw_133_module_data_out[4] ,
    \sw_133_module_data_out[3] ,
    \sw_133_module_data_out[2] ,
    \sw_133_module_data_out[1] ,
    \sw_133_module_data_out[0] }));
 scanchain scanchain_134 (.clk_in(sw_133_clk_out),
    .clk_out(sw_134_clk_out),
    .data_in(sw_133_data_out),
    .data_out(sw_134_data_out),
    .latch_enable_in(sw_133_latch_out),
    .latch_enable_out(sw_134_latch_out),
    .scan_select_in(sw_133_scan_out),
    .scan_select_out(sw_134_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_134_module_data_in[7] ,
    \sw_134_module_data_in[6] ,
    \sw_134_module_data_in[5] ,
    \sw_134_module_data_in[4] ,
    \sw_134_module_data_in[3] ,
    \sw_134_module_data_in[2] ,
    \sw_134_module_data_in[1] ,
    \sw_134_module_data_in[0] }),
    .module_data_out({\sw_134_module_data_out[7] ,
    \sw_134_module_data_out[6] ,
    \sw_134_module_data_out[5] ,
    \sw_134_module_data_out[4] ,
    \sw_134_module_data_out[3] ,
    \sw_134_module_data_out[2] ,
    \sw_134_module_data_out[1] ,
    \sw_134_module_data_out[0] }));
 scanchain scanchain_135 (.clk_in(sw_134_clk_out),
    .clk_out(sw_135_clk_out),
    .data_in(sw_134_data_out),
    .data_out(sw_135_data_out),
    .latch_enable_in(sw_134_latch_out),
    .latch_enable_out(sw_135_latch_out),
    .scan_select_in(sw_134_scan_out),
    .scan_select_out(sw_135_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_135_module_data_in[7] ,
    \sw_135_module_data_in[6] ,
    \sw_135_module_data_in[5] ,
    \sw_135_module_data_in[4] ,
    \sw_135_module_data_in[3] ,
    \sw_135_module_data_in[2] ,
    \sw_135_module_data_in[1] ,
    \sw_135_module_data_in[0] }),
    .module_data_out({\sw_135_module_data_out[7] ,
    \sw_135_module_data_out[6] ,
    \sw_135_module_data_out[5] ,
    \sw_135_module_data_out[4] ,
    \sw_135_module_data_out[3] ,
    \sw_135_module_data_out[2] ,
    \sw_135_module_data_out[1] ,
    \sw_135_module_data_out[0] }));
 scanchain scanchain_136 (.clk_in(sw_135_clk_out),
    .clk_out(sw_136_clk_out),
    .data_in(sw_135_data_out),
    .data_out(sw_136_data_out),
    .latch_enable_in(sw_135_latch_out),
    .latch_enable_out(sw_136_latch_out),
    .scan_select_in(sw_135_scan_out),
    .scan_select_out(sw_136_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_136_module_data_in[7] ,
    \sw_136_module_data_in[6] ,
    \sw_136_module_data_in[5] ,
    \sw_136_module_data_in[4] ,
    \sw_136_module_data_in[3] ,
    \sw_136_module_data_in[2] ,
    \sw_136_module_data_in[1] ,
    \sw_136_module_data_in[0] }),
    .module_data_out({\sw_136_module_data_out[7] ,
    \sw_136_module_data_out[6] ,
    \sw_136_module_data_out[5] ,
    \sw_136_module_data_out[4] ,
    \sw_136_module_data_out[3] ,
    \sw_136_module_data_out[2] ,
    \sw_136_module_data_out[1] ,
    \sw_136_module_data_out[0] }));
 scanchain scanchain_137 (.clk_in(sw_136_clk_out),
    .clk_out(sw_137_clk_out),
    .data_in(sw_136_data_out),
    .data_out(sw_137_data_out),
    .latch_enable_in(sw_136_latch_out),
    .latch_enable_out(sw_137_latch_out),
    .scan_select_in(sw_136_scan_out),
    .scan_select_out(sw_137_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_137_module_data_in[7] ,
    \sw_137_module_data_in[6] ,
    \sw_137_module_data_in[5] ,
    \sw_137_module_data_in[4] ,
    \sw_137_module_data_in[3] ,
    \sw_137_module_data_in[2] ,
    \sw_137_module_data_in[1] ,
    \sw_137_module_data_in[0] }),
    .module_data_out({\sw_137_module_data_out[7] ,
    \sw_137_module_data_out[6] ,
    \sw_137_module_data_out[5] ,
    \sw_137_module_data_out[4] ,
    \sw_137_module_data_out[3] ,
    \sw_137_module_data_out[2] ,
    \sw_137_module_data_out[1] ,
    \sw_137_module_data_out[0] }));
 scanchain scanchain_138 (.clk_in(sw_137_clk_out),
    .clk_out(sw_138_clk_out),
    .data_in(sw_137_data_out),
    .data_out(sw_138_data_out),
    .latch_enable_in(sw_137_latch_out),
    .latch_enable_out(sw_138_latch_out),
    .scan_select_in(sw_137_scan_out),
    .scan_select_out(sw_138_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_138_module_data_in[7] ,
    \sw_138_module_data_in[6] ,
    \sw_138_module_data_in[5] ,
    \sw_138_module_data_in[4] ,
    \sw_138_module_data_in[3] ,
    \sw_138_module_data_in[2] ,
    \sw_138_module_data_in[1] ,
    \sw_138_module_data_in[0] }),
    .module_data_out({\sw_138_module_data_out[7] ,
    \sw_138_module_data_out[6] ,
    \sw_138_module_data_out[5] ,
    \sw_138_module_data_out[4] ,
    \sw_138_module_data_out[3] ,
    \sw_138_module_data_out[2] ,
    \sw_138_module_data_out[1] ,
    \sw_138_module_data_out[0] }));
 scanchain scanchain_139 (.clk_in(sw_138_clk_out),
    .clk_out(sw_139_clk_out),
    .data_in(sw_138_data_out),
    .data_out(sw_139_data_out),
    .latch_enable_in(sw_138_latch_out),
    .latch_enable_out(sw_139_latch_out),
    .scan_select_in(sw_138_scan_out),
    .scan_select_out(sw_139_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_139_module_data_in[7] ,
    \sw_139_module_data_in[6] ,
    \sw_139_module_data_in[5] ,
    \sw_139_module_data_in[4] ,
    \sw_139_module_data_in[3] ,
    \sw_139_module_data_in[2] ,
    \sw_139_module_data_in[1] ,
    \sw_139_module_data_in[0] }),
    .module_data_out({\sw_139_module_data_out[7] ,
    \sw_139_module_data_out[6] ,
    \sw_139_module_data_out[5] ,
    \sw_139_module_data_out[4] ,
    \sw_139_module_data_out[3] ,
    \sw_139_module_data_out[2] ,
    \sw_139_module_data_out[1] ,
    \sw_139_module_data_out[0] }));
 scanchain scanchain_140 (.clk_in(sw_139_clk_out),
    .clk_out(sw_140_clk_out),
    .data_in(sw_139_data_out),
    .data_out(sw_140_data_out),
    .latch_enable_in(sw_139_latch_out),
    .latch_enable_out(sw_140_latch_out),
    .scan_select_in(sw_139_scan_out),
    .scan_select_out(sw_140_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_140_module_data_in[7] ,
    \sw_140_module_data_in[6] ,
    \sw_140_module_data_in[5] ,
    \sw_140_module_data_in[4] ,
    \sw_140_module_data_in[3] ,
    \sw_140_module_data_in[2] ,
    \sw_140_module_data_in[1] ,
    \sw_140_module_data_in[0] }),
    .module_data_out({\sw_140_module_data_out[7] ,
    \sw_140_module_data_out[6] ,
    \sw_140_module_data_out[5] ,
    \sw_140_module_data_out[4] ,
    \sw_140_module_data_out[3] ,
    \sw_140_module_data_out[2] ,
    \sw_140_module_data_out[1] ,
    \sw_140_module_data_out[0] }));
 scanchain scanchain_141 (.clk_in(sw_140_clk_out),
    .clk_out(sw_141_clk_out),
    .data_in(sw_140_data_out),
    .data_out(sw_141_data_out),
    .latch_enable_in(sw_140_latch_out),
    .latch_enable_out(sw_141_latch_out),
    .scan_select_in(sw_140_scan_out),
    .scan_select_out(sw_141_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_141_module_data_in[7] ,
    \sw_141_module_data_in[6] ,
    \sw_141_module_data_in[5] ,
    \sw_141_module_data_in[4] ,
    \sw_141_module_data_in[3] ,
    \sw_141_module_data_in[2] ,
    \sw_141_module_data_in[1] ,
    \sw_141_module_data_in[0] }),
    .module_data_out({\sw_141_module_data_out[7] ,
    \sw_141_module_data_out[6] ,
    \sw_141_module_data_out[5] ,
    \sw_141_module_data_out[4] ,
    \sw_141_module_data_out[3] ,
    \sw_141_module_data_out[2] ,
    \sw_141_module_data_out[1] ,
    \sw_141_module_data_out[0] }));
 scanchain scanchain_142 (.clk_in(sw_141_clk_out),
    .clk_out(sw_142_clk_out),
    .data_in(sw_141_data_out),
    .data_out(sw_142_data_out),
    .latch_enable_in(sw_141_latch_out),
    .latch_enable_out(sw_142_latch_out),
    .scan_select_in(sw_141_scan_out),
    .scan_select_out(sw_142_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_142_module_data_in[7] ,
    \sw_142_module_data_in[6] ,
    \sw_142_module_data_in[5] ,
    \sw_142_module_data_in[4] ,
    \sw_142_module_data_in[3] ,
    \sw_142_module_data_in[2] ,
    \sw_142_module_data_in[1] ,
    \sw_142_module_data_in[0] }),
    .module_data_out({\sw_142_module_data_out[7] ,
    \sw_142_module_data_out[6] ,
    \sw_142_module_data_out[5] ,
    \sw_142_module_data_out[4] ,
    \sw_142_module_data_out[3] ,
    \sw_142_module_data_out[2] ,
    \sw_142_module_data_out[1] ,
    \sw_142_module_data_out[0] }));
 scanchain scanchain_143 (.clk_in(sw_142_clk_out),
    .clk_out(sw_143_clk_out),
    .data_in(sw_142_data_out),
    .data_out(sw_143_data_out),
    .latch_enable_in(sw_142_latch_out),
    .latch_enable_out(sw_143_latch_out),
    .scan_select_in(sw_142_scan_out),
    .scan_select_out(sw_143_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_143_module_data_in[7] ,
    \sw_143_module_data_in[6] ,
    \sw_143_module_data_in[5] ,
    \sw_143_module_data_in[4] ,
    \sw_143_module_data_in[3] ,
    \sw_143_module_data_in[2] ,
    \sw_143_module_data_in[1] ,
    \sw_143_module_data_in[0] }),
    .module_data_out({\sw_143_module_data_out[7] ,
    \sw_143_module_data_out[6] ,
    \sw_143_module_data_out[5] ,
    \sw_143_module_data_out[4] ,
    \sw_143_module_data_out[3] ,
    \sw_143_module_data_out[2] ,
    \sw_143_module_data_out[1] ,
    \sw_143_module_data_out[0] }));
 scanchain scanchain_144 (.clk_in(sw_143_clk_out),
    .clk_out(sw_144_clk_out),
    .data_in(sw_143_data_out),
    .data_out(sw_144_data_out),
    .latch_enable_in(sw_143_latch_out),
    .latch_enable_out(sw_144_latch_out),
    .scan_select_in(sw_143_scan_out),
    .scan_select_out(sw_144_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_144_module_data_in[7] ,
    \sw_144_module_data_in[6] ,
    \sw_144_module_data_in[5] ,
    \sw_144_module_data_in[4] ,
    \sw_144_module_data_in[3] ,
    \sw_144_module_data_in[2] ,
    \sw_144_module_data_in[1] ,
    \sw_144_module_data_in[0] }),
    .module_data_out({\sw_144_module_data_out[7] ,
    \sw_144_module_data_out[6] ,
    \sw_144_module_data_out[5] ,
    \sw_144_module_data_out[4] ,
    \sw_144_module_data_out[3] ,
    \sw_144_module_data_out[2] ,
    \sw_144_module_data_out[1] ,
    \sw_144_module_data_out[0] }));
 scanchain scanchain_145 (.clk_in(sw_144_clk_out),
    .clk_out(sw_145_clk_out),
    .data_in(sw_144_data_out),
    .data_out(sw_145_data_out),
    .latch_enable_in(sw_144_latch_out),
    .latch_enable_out(sw_145_latch_out),
    .scan_select_in(sw_144_scan_out),
    .scan_select_out(sw_145_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_145_module_data_in[7] ,
    \sw_145_module_data_in[6] ,
    \sw_145_module_data_in[5] ,
    \sw_145_module_data_in[4] ,
    \sw_145_module_data_in[3] ,
    \sw_145_module_data_in[2] ,
    \sw_145_module_data_in[1] ,
    \sw_145_module_data_in[0] }),
    .module_data_out({\sw_145_module_data_out[7] ,
    \sw_145_module_data_out[6] ,
    \sw_145_module_data_out[5] ,
    \sw_145_module_data_out[4] ,
    \sw_145_module_data_out[3] ,
    \sw_145_module_data_out[2] ,
    \sw_145_module_data_out[1] ,
    \sw_145_module_data_out[0] }));
 scanchain scanchain_146 (.clk_in(sw_145_clk_out),
    .clk_out(sw_146_clk_out),
    .data_in(sw_145_data_out),
    .data_out(sw_146_data_out),
    .latch_enable_in(sw_145_latch_out),
    .latch_enable_out(sw_146_latch_out),
    .scan_select_in(sw_145_scan_out),
    .scan_select_out(sw_146_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_146_module_data_in[7] ,
    \sw_146_module_data_in[6] ,
    \sw_146_module_data_in[5] ,
    \sw_146_module_data_in[4] ,
    \sw_146_module_data_in[3] ,
    \sw_146_module_data_in[2] ,
    \sw_146_module_data_in[1] ,
    \sw_146_module_data_in[0] }),
    .module_data_out({\sw_146_module_data_out[7] ,
    \sw_146_module_data_out[6] ,
    \sw_146_module_data_out[5] ,
    \sw_146_module_data_out[4] ,
    \sw_146_module_data_out[3] ,
    \sw_146_module_data_out[2] ,
    \sw_146_module_data_out[1] ,
    \sw_146_module_data_out[0] }));
 scanchain scanchain_147 (.clk_in(sw_146_clk_out),
    .clk_out(sw_147_clk_out),
    .data_in(sw_146_data_out),
    .data_out(sw_147_data_out),
    .latch_enable_in(sw_146_latch_out),
    .latch_enable_out(sw_147_latch_out),
    .scan_select_in(sw_146_scan_out),
    .scan_select_out(sw_147_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_147_module_data_in[7] ,
    \sw_147_module_data_in[6] ,
    \sw_147_module_data_in[5] ,
    \sw_147_module_data_in[4] ,
    \sw_147_module_data_in[3] ,
    \sw_147_module_data_in[2] ,
    \sw_147_module_data_in[1] ,
    \sw_147_module_data_in[0] }),
    .module_data_out({\sw_147_module_data_out[7] ,
    \sw_147_module_data_out[6] ,
    \sw_147_module_data_out[5] ,
    \sw_147_module_data_out[4] ,
    \sw_147_module_data_out[3] ,
    \sw_147_module_data_out[2] ,
    \sw_147_module_data_out[1] ,
    \sw_147_module_data_out[0] }));
 scanchain scanchain_148 (.clk_in(sw_147_clk_out),
    .clk_out(sw_148_clk_out),
    .data_in(sw_147_data_out),
    .data_out(sw_148_data_out),
    .latch_enable_in(sw_147_latch_out),
    .latch_enable_out(sw_148_latch_out),
    .scan_select_in(sw_147_scan_out),
    .scan_select_out(sw_148_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_148_module_data_in[7] ,
    \sw_148_module_data_in[6] ,
    \sw_148_module_data_in[5] ,
    \sw_148_module_data_in[4] ,
    \sw_148_module_data_in[3] ,
    \sw_148_module_data_in[2] ,
    \sw_148_module_data_in[1] ,
    \sw_148_module_data_in[0] }),
    .module_data_out({\sw_148_module_data_out[7] ,
    \sw_148_module_data_out[6] ,
    \sw_148_module_data_out[5] ,
    \sw_148_module_data_out[4] ,
    \sw_148_module_data_out[3] ,
    \sw_148_module_data_out[2] ,
    \sw_148_module_data_out[1] ,
    \sw_148_module_data_out[0] }));
 scanchain scanchain_149 (.clk_in(sw_148_clk_out),
    .clk_out(sw_149_clk_out),
    .data_in(sw_148_data_out),
    .data_out(sw_149_data_out),
    .latch_enable_in(sw_148_latch_out),
    .latch_enable_out(sw_149_latch_out),
    .scan_select_in(sw_148_scan_out),
    .scan_select_out(sw_149_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_149_module_data_in[7] ,
    \sw_149_module_data_in[6] ,
    \sw_149_module_data_in[5] ,
    \sw_149_module_data_in[4] ,
    \sw_149_module_data_in[3] ,
    \sw_149_module_data_in[2] ,
    \sw_149_module_data_in[1] ,
    \sw_149_module_data_in[0] }),
    .module_data_out({\sw_149_module_data_out[7] ,
    \sw_149_module_data_out[6] ,
    \sw_149_module_data_out[5] ,
    \sw_149_module_data_out[4] ,
    \sw_149_module_data_out[3] ,
    \sw_149_module_data_out[2] ,
    \sw_149_module_data_out[1] ,
    \sw_149_module_data_out[0] }));
 scanchain scanchain_150 (.clk_in(sw_149_clk_out),
    .clk_out(sw_150_clk_out),
    .data_in(sw_149_data_out),
    .data_out(sw_150_data_out),
    .latch_enable_in(sw_149_latch_out),
    .latch_enable_out(sw_150_latch_out),
    .scan_select_in(sw_149_scan_out),
    .scan_select_out(sw_150_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_150_module_data_in[7] ,
    \sw_150_module_data_in[6] ,
    \sw_150_module_data_in[5] ,
    \sw_150_module_data_in[4] ,
    \sw_150_module_data_in[3] ,
    \sw_150_module_data_in[2] ,
    \sw_150_module_data_in[1] ,
    \sw_150_module_data_in[0] }),
    .module_data_out({\sw_150_module_data_out[7] ,
    \sw_150_module_data_out[6] ,
    \sw_150_module_data_out[5] ,
    \sw_150_module_data_out[4] ,
    \sw_150_module_data_out[3] ,
    \sw_150_module_data_out[2] ,
    \sw_150_module_data_out[1] ,
    \sw_150_module_data_out[0] }));
 scanchain scanchain_151 (.clk_in(sw_150_clk_out),
    .clk_out(sw_151_clk_out),
    .data_in(sw_150_data_out),
    .data_out(sw_151_data_out),
    .latch_enable_in(sw_150_latch_out),
    .latch_enable_out(sw_151_latch_out),
    .scan_select_in(sw_150_scan_out),
    .scan_select_out(sw_151_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_151_module_data_in[7] ,
    \sw_151_module_data_in[6] ,
    \sw_151_module_data_in[5] ,
    \sw_151_module_data_in[4] ,
    \sw_151_module_data_in[3] ,
    \sw_151_module_data_in[2] ,
    \sw_151_module_data_in[1] ,
    \sw_151_module_data_in[0] }),
    .module_data_out({\sw_151_module_data_out[7] ,
    \sw_151_module_data_out[6] ,
    \sw_151_module_data_out[5] ,
    \sw_151_module_data_out[4] ,
    \sw_151_module_data_out[3] ,
    \sw_151_module_data_out[2] ,
    \sw_151_module_data_out[1] ,
    \sw_151_module_data_out[0] }));
 scanchain scanchain_152 (.clk_in(sw_151_clk_out),
    .clk_out(sw_152_clk_out),
    .data_in(sw_151_data_out),
    .data_out(sw_152_data_out),
    .latch_enable_in(sw_151_latch_out),
    .latch_enable_out(sw_152_latch_out),
    .scan_select_in(sw_151_scan_out),
    .scan_select_out(sw_152_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_152_module_data_in[7] ,
    \sw_152_module_data_in[6] ,
    \sw_152_module_data_in[5] ,
    \sw_152_module_data_in[4] ,
    \sw_152_module_data_in[3] ,
    \sw_152_module_data_in[2] ,
    \sw_152_module_data_in[1] ,
    \sw_152_module_data_in[0] }),
    .module_data_out({\sw_152_module_data_out[7] ,
    \sw_152_module_data_out[6] ,
    \sw_152_module_data_out[5] ,
    \sw_152_module_data_out[4] ,
    \sw_152_module_data_out[3] ,
    \sw_152_module_data_out[2] ,
    \sw_152_module_data_out[1] ,
    \sw_152_module_data_out[0] }));
 scanchain scanchain_153 (.clk_in(sw_152_clk_out),
    .clk_out(sw_153_clk_out),
    .data_in(sw_152_data_out),
    .data_out(sw_153_data_out),
    .latch_enable_in(sw_152_latch_out),
    .latch_enable_out(sw_153_latch_out),
    .scan_select_in(sw_152_scan_out),
    .scan_select_out(sw_153_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_153_module_data_in[7] ,
    \sw_153_module_data_in[6] ,
    \sw_153_module_data_in[5] ,
    \sw_153_module_data_in[4] ,
    \sw_153_module_data_in[3] ,
    \sw_153_module_data_in[2] ,
    \sw_153_module_data_in[1] ,
    \sw_153_module_data_in[0] }),
    .module_data_out({\sw_153_module_data_out[7] ,
    \sw_153_module_data_out[6] ,
    \sw_153_module_data_out[5] ,
    \sw_153_module_data_out[4] ,
    \sw_153_module_data_out[3] ,
    \sw_153_module_data_out[2] ,
    \sw_153_module_data_out[1] ,
    \sw_153_module_data_out[0] }));
 scanchain scanchain_154 (.clk_in(sw_153_clk_out),
    .clk_out(sw_154_clk_out),
    .data_in(sw_153_data_out),
    .data_out(sw_154_data_out),
    .latch_enable_in(sw_153_latch_out),
    .latch_enable_out(sw_154_latch_out),
    .scan_select_in(sw_153_scan_out),
    .scan_select_out(sw_154_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_154_module_data_in[7] ,
    \sw_154_module_data_in[6] ,
    \sw_154_module_data_in[5] ,
    \sw_154_module_data_in[4] ,
    \sw_154_module_data_in[3] ,
    \sw_154_module_data_in[2] ,
    \sw_154_module_data_in[1] ,
    \sw_154_module_data_in[0] }),
    .module_data_out({\sw_154_module_data_out[7] ,
    \sw_154_module_data_out[6] ,
    \sw_154_module_data_out[5] ,
    \sw_154_module_data_out[4] ,
    \sw_154_module_data_out[3] ,
    \sw_154_module_data_out[2] ,
    \sw_154_module_data_out[1] ,
    \sw_154_module_data_out[0] }));
 scanchain scanchain_155 (.clk_in(sw_154_clk_out),
    .clk_out(sw_155_clk_out),
    .data_in(sw_154_data_out),
    .data_out(sw_155_data_out),
    .latch_enable_in(sw_154_latch_out),
    .latch_enable_out(sw_155_latch_out),
    .scan_select_in(sw_154_scan_out),
    .scan_select_out(sw_155_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_155_module_data_in[7] ,
    \sw_155_module_data_in[6] ,
    \sw_155_module_data_in[5] ,
    \sw_155_module_data_in[4] ,
    \sw_155_module_data_in[3] ,
    \sw_155_module_data_in[2] ,
    \sw_155_module_data_in[1] ,
    \sw_155_module_data_in[0] }),
    .module_data_out({\sw_155_module_data_out[7] ,
    \sw_155_module_data_out[6] ,
    \sw_155_module_data_out[5] ,
    \sw_155_module_data_out[4] ,
    \sw_155_module_data_out[3] ,
    \sw_155_module_data_out[2] ,
    \sw_155_module_data_out[1] ,
    \sw_155_module_data_out[0] }));
 scanchain scanchain_156 (.clk_in(sw_155_clk_out),
    .clk_out(sw_156_clk_out),
    .data_in(sw_155_data_out),
    .data_out(sw_156_data_out),
    .latch_enable_in(sw_155_latch_out),
    .latch_enable_out(sw_156_latch_out),
    .scan_select_in(sw_155_scan_out),
    .scan_select_out(sw_156_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_156_module_data_in[7] ,
    \sw_156_module_data_in[6] ,
    \sw_156_module_data_in[5] ,
    \sw_156_module_data_in[4] ,
    \sw_156_module_data_in[3] ,
    \sw_156_module_data_in[2] ,
    \sw_156_module_data_in[1] ,
    \sw_156_module_data_in[0] }),
    .module_data_out({\sw_156_module_data_out[7] ,
    \sw_156_module_data_out[6] ,
    \sw_156_module_data_out[5] ,
    \sw_156_module_data_out[4] ,
    \sw_156_module_data_out[3] ,
    \sw_156_module_data_out[2] ,
    \sw_156_module_data_out[1] ,
    \sw_156_module_data_out[0] }));
 scanchain scanchain_157 (.clk_in(sw_156_clk_out),
    .clk_out(sw_157_clk_out),
    .data_in(sw_156_data_out),
    .data_out(sw_157_data_out),
    .latch_enable_in(sw_156_latch_out),
    .latch_enable_out(sw_157_latch_out),
    .scan_select_in(sw_156_scan_out),
    .scan_select_out(sw_157_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_157_module_data_in[7] ,
    \sw_157_module_data_in[6] ,
    \sw_157_module_data_in[5] ,
    \sw_157_module_data_in[4] ,
    \sw_157_module_data_in[3] ,
    \sw_157_module_data_in[2] ,
    \sw_157_module_data_in[1] ,
    \sw_157_module_data_in[0] }),
    .module_data_out({\sw_157_module_data_out[7] ,
    \sw_157_module_data_out[6] ,
    \sw_157_module_data_out[5] ,
    \sw_157_module_data_out[4] ,
    \sw_157_module_data_out[3] ,
    \sw_157_module_data_out[2] ,
    \sw_157_module_data_out[1] ,
    \sw_157_module_data_out[0] }));
 scanchain scanchain_158 (.clk_in(sw_157_clk_out),
    .clk_out(sw_158_clk_out),
    .data_in(sw_157_data_out),
    .data_out(sw_158_data_out),
    .latch_enable_in(sw_157_latch_out),
    .latch_enable_out(sw_158_latch_out),
    .scan_select_in(sw_157_scan_out),
    .scan_select_out(sw_158_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_158_module_data_in[7] ,
    \sw_158_module_data_in[6] ,
    \sw_158_module_data_in[5] ,
    \sw_158_module_data_in[4] ,
    \sw_158_module_data_in[3] ,
    \sw_158_module_data_in[2] ,
    \sw_158_module_data_in[1] ,
    \sw_158_module_data_in[0] }),
    .module_data_out({\sw_158_module_data_out[7] ,
    \sw_158_module_data_out[6] ,
    \sw_158_module_data_out[5] ,
    \sw_158_module_data_out[4] ,
    \sw_158_module_data_out[3] ,
    \sw_158_module_data_out[2] ,
    \sw_158_module_data_out[1] ,
    \sw_158_module_data_out[0] }));
 scanchain scanchain_159 (.clk_in(sw_158_clk_out),
    .clk_out(sw_159_clk_out),
    .data_in(sw_158_data_out),
    .data_out(sw_159_data_out),
    .latch_enable_in(sw_158_latch_out),
    .latch_enable_out(sw_159_latch_out),
    .scan_select_in(sw_158_scan_out),
    .scan_select_out(sw_159_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_159_module_data_in[7] ,
    \sw_159_module_data_in[6] ,
    \sw_159_module_data_in[5] ,
    \sw_159_module_data_in[4] ,
    \sw_159_module_data_in[3] ,
    \sw_159_module_data_in[2] ,
    \sw_159_module_data_in[1] ,
    \sw_159_module_data_in[0] }),
    .module_data_out({\sw_159_module_data_out[7] ,
    \sw_159_module_data_out[6] ,
    \sw_159_module_data_out[5] ,
    \sw_159_module_data_out[4] ,
    \sw_159_module_data_out[3] ,
    \sw_159_module_data_out[2] ,
    \sw_159_module_data_out[1] ,
    \sw_159_module_data_out[0] }));
 scanchain scanchain_160 (.clk_in(sw_159_clk_out),
    .clk_out(sw_160_clk_out),
    .data_in(sw_159_data_out),
    .data_out(sw_160_data_out),
    .latch_enable_in(sw_159_latch_out),
    .latch_enable_out(sw_160_latch_out),
    .scan_select_in(sw_159_scan_out),
    .scan_select_out(sw_160_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_160_module_data_in[7] ,
    \sw_160_module_data_in[6] ,
    \sw_160_module_data_in[5] ,
    \sw_160_module_data_in[4] ,
    \sw_160_module_data_in[3] ,
    \sw_160_module_data_in[2] ,
    \sw_160_module_data_in[1] ,
    \sw_160_module_data_in[0] }),
    .module_data_out({\sw_160_module_data_out[7] ,
    \sw_160_module_data_out[6] ,
    \sw_160_module_data_out[5] ,
    \sw_160_module_data_out[4] ,
    \sw_160_module_data_out[3] ,
    \sw_160_module_data_out[2] ,
    \sw_160_module_data_out[1] ,
    \sw_160_module_data_out[0] }));
 scanchain scanchain_161 (.clk_in(sw_160_clk_out),
    .clk_out(sw_161_clk_out),
    .data_in(sw_160_data_out),
    .data_out(sw_161_data_out),
    .latch_enable_in(sw_160_latch_out),
    .latch_enable_out(sw_161_latch_out),
    .scan_select_in(sw_160_scan_out),
    .scan_select_out(sw_161_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_161_module_data_in[7] ,
    \sw_161_module_data_in[6] ,
    \sw_161_module_data_in[5] ,
    \sw_161_module_data_in[4] ,
    \sw_161_module_data_in[3] ,
    \sw_161_module_data_in[2] ,
    \sw_161_module_data_in[1] ,
    \sw_161_module_data_in[0] }),
    .module_data_out({\sw_161_module_data_out[7] ,
    \sw_161_module_data_out[6] ,
    \sw_161_module_data_out[5] ,
    \sw_161_module_data_out[4] ,
    \sw_161_module_data_out[3] ,
    \sw_161_module_data_out[2] ,
    \sw_161_module_data_out[1] ,
    \sw_161_module_data_out[0] }));
 scanchain scanchain_162 (.clk_in(sw_161_clk_out),
    .clk_out(sw_162_clk_out),
    .data_in(sw_161_data_out),
    .data_out(sw_162_data_out),
    .latch_enable_in(sw_161_latch_out),
    .latch_enable_out(sw_162_latch_out),
    .scan_select_in(sw_161_scan_out),
    .scan_select_out(sw_162_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_162_module_data_in[7] ,
    \sw_162_module_data_in[6] ,
    \sw_162_module_data_in[5] ,
    \sw_162_module_data_in[4] ,
    \sw_162_module_data_in[3] ,
    \sw_162_module_data_in[2] ,
    \sw_162_module_data_in[1] ,
    \sw_162_module_data_in[0] }),
    .module_data_out({\sw_162_module_data_out[7] ,
    \sw_162_module_data_out[6] ,
    \sw_162_module_data_out[5] ,
    \sw_162_module_data_out[4] ,
    \sw_162_module_data_out[3] ,
    \sw_162_module_data_out[2] ,
    \sw_162_module_data_out[1] ,
    \sw_162_module_data_out[0] }));
 scanchain scanchain_163 (.clk_in(sw_162_clk_out),
    .clk_out(sw_163_clk_out),
    .data_in(sw_162_data_out),
    .data_out(sw_163_data_out),
    .latch_enable_in(sw_162_latch_out),
    .latch_enable_out(sw_163_latch_out),
    .scan_select_in(sw_162_scan_out),
    .scan_select_out(sw_163_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_163_module_data_in[7] ,
    \sw_163_module_data_in[6] ,
    \sw_163_module_data_in[5] ,
    \sw_163_module_data_in[4] ,
    \sw_163_module_data_in[3] ,
    \sw_163_module_data_in[2] ,
    \sw_163_module_data_in[1] ,
    \sw_163_module_data_in[0] }),
    .module_data_out({\sw_163_module_data_out[7] ,
    \sw_163_module_data_out[6] ,
    \sw_163_module_data_out[5] ,
    \sw_163_module_data_out[4] ,
    \sw_163_module_data_out[3] ,
    \sw_163_module_data_out[2] ,
    \sw_163_module_data_out[1] ,
    \sw_163_module_data_out[0] }));
 scanchain scanchain_164 (.clk_in(sw_163_clk_out),
    .clk_out(sw_164_clk_out),
    .data_in(sw_163_data_out),
    .data_out(sw_164_data_out),
    .latch_enable_in(sw_163_latch_out),
    .latch_enable_out(sw_164_latch_out),
    .scan_select_in(sw_163_scan_out),
    .scan_select_out(sw_164_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_164_module_data_in[7] ,
    \sw_164_module_data_in[6] ,
    \sw_164_module_data_in[5] ,
    \sw_164_module_data_in[4] ,
    \sw_164_module_data_in[3] ,
    \sw_164_module_data_in[2] ,
    \sw_164_module_data_in[1] ,
    \sw_164_module_data_in[0] }),
    .module_data_out({\sw_164_module_data_out[7] ,
    \sw_164_module_data_out[6] ,
    \sw_164_module_data_out[5] ,
    \sw_164_module_data_out[4] ,
    \sw_164_module_data_out[3] ,
    \sw_164_module_data_out[2] ,
    \sw_164_module_data_out[1] ,
    \sw_164_module_data_out[0] }));
 scanchain scanchain_165 (.clk_in(sw_164_clk_out),
    .clk_out(sw_165_clk_out),
    .data_in(sw_164_data_out),
    .data_out(sw_165_data_out),
    .latch_enable_in(sw_164_latch_out),
    .latch_enable_out(sw_165_latch_out),
    .scan_select_in(sw_164_scan_out),
    .scan_select_out(sw_165_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_165_module_data_in[7] ,
    \sw_165_module_data_in[6] ,
    \sw_165_module_data_in[5] ,
    \sw_165_module_data_in[4] ,
    \sw_165_module_data_in[3] ,
    \sw_165_module_data_in[2] ,
    \sw_165_module_data_in[1] ,
    \sw_165_module_data_in[0] }),
    .module_data_out({\sw_165_module_data_out[7] ,
    \sw_165_module_data_out[6] ,
    \sw_165_module_data_out[5] ,
    \sw_165_module_data_out[4] ,
    \sw_165_module_data_out[3] ,
    \sw_165_module_data_out[2] ,
    \sw_165_module_data_out[1] ,
    \sw_165_module_data_out[0] }));
 scanchain scanchain_166 (.clk_in(sw_165_clk_out),
    .clk_out(sw_166_clk_out),
    .data_in(sw_165_data_out),
    .data_out(sw_166_data_out),
    .latch_enable_in(sw_165_latch_out),
    .latch_enable_out(sw_166_latch_out),
    .scan_select_in(sw_165_scan_out),
    .scan_select_out(sw_166_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_166_module_data_in[7] ,
    \sw_166_module_data_in[6] ,
    \sw_166_module_data_in[5] ,
    \sw_166_module_data_in[4] ,
    \sw_166_module_data_in[3] ,
    \sw_166_module_data_in[2] ,
    \sw_166_module_data_in[1] ,
    \sw_166_module_data_in[0] }),
    .module_data_out({\sw_166_module_data_out[7] ,
    \sw_166_module_data_out[6] ,
    \sw_166_module_data_out[5] ,
    \sw_166_module_data_out[4] ,
    \sw_166_module_data_out[3] ,
    \sw_166_module_data_out[2] ,
    \sw_166_module_data_out[1] ,
    \sw_166_module_data_out[0] }));
 scanchain scanchain_167 (.clk_in(sw_166_clk_out),
    .clk_out(sw_167_clk_out),
    .data_in(sw_166_data_out),
    .data_out(sw_167_data_out),
    .latch_enable_in(sw_166_latch_out),
    .latch_enable_out(sw_167_latch_out),
    .scan_select_in(sw_166_scan_out),
    .scan_select_out(sw_167_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_167_module_data_in[7] ,
    \sw_167_module_data_in[6] ,
    \sw_167_module_data_in[5] ,
    \sw_167_module_data_in[4] ,
    \sw_167_module_data_in[3] ,
    \sw_167_module_data_in[2] ,
    \sw_167_module_data_in[1] ,
    \sw_167_module_data_in[0] }),
    .module_data_out({\sw_167_module_data_out[7] ,
    \sw_167_module_data_out[6] ,
    \sw_167_module_data_out[5] ,
    \sw_167_module_data_out[4] ,
    \sw_167_module_data_out[3] ,
    \sw_167_module_data_out[2] ,
    \sw_167_module_data_out[1] ,
    \sw_167_module_data_out[0] }));
 scanchain scanchain_168 (.clk_in(sw_167_clk_out),
    .clk_out(sw_168_clk_out),
    .data_in(sw_167_data_out),
    .data_out(sw_168_data_out),
    .latch_enable_in(sw_167_latch_out),
    .latch_enable_out(sw_168_latch_out),
    .scan_select_in(sw_167_scan_out),
    .scan_select_out(sw_168_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_168_module_data_in[7] ,
    \sw_168_module_data_in[6] ,
    \sw_168_module_data_in[5] ,
    \sw_168_module_data_in[4] ,
    \sw_168_module_data_in[3] ,
    \sw_168_module_data_in[2] ,
    \sw_168_module_data_in[1] ,
    \sw_168_module_data_in[0] }),
    .module_data_out({\sw_168_module_data_out[7] ,
    \sw_168_module_data_out[6] ,
    \sw_168_module_data_out[5] ,
    \sw_168_module_data_out[4] ,
    \sw_168_module_data_out[3] ,
    \sw_168_module_data_out[2] ,
    \sw_168_module_data_out[1] ,
    \sw_168_module_data_out[0] }));
 scanchain scanchain_169 (.clk_in(sw_168_clk_out),
    .clk_out(sw_169_clk_out),
    .data_in(sw_168_data_out),
    .data_out(sw_169_data_out),
    .latch_enable_in(sw_168_latch_out),
    .latch_enable_out(sw_169_latch_out),
    .scan_select_in(sw_168_scan_out),
    .scan_select_out(sw_169_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_169_module_data_in[7] ,
    \sw_169_module_data_in[6] ,
    \sw_169_module_data_in[5] ,
    \sw_169_module_data_in[4] ,
    \sw_169_module_data_in[3] ,
    \sw_169_module_data_in[2] ,
    \sw_169_module_data_in[1] ,
    \sw_169_module_data_in[0] }),
    .module_data_out({\sw_169_module_data_out[7] ,
    \sw_169_module_data_out[6] ,
    \sw_169_module_data_out[5] ,
    \sw_169_module_data_out[4] ,
    \sw_169_module_data_out[3] ,
    \sw_169_module_data_out[2] ,
    \sw_169_module_data_out[1] ,
    \sw_169_module_data_out[0] }));
 scanchain scanchain_170 (.clk_in(sw_169_clk_out),
    .clk_out(sw_170_clk_out),
    .data_in(sw_169_data_out),
    .data_out(sw_170_data_out),
    .latch_enable_in(sw_169_latch_out),
    .latch_enable_out(sw_170_latch_out),
    .scan_select_in(sw_169_scan_out),
    .scan_select_out(sw_170_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_170_module_data_in[7] ,
    \sw_170_module_data_in[6] ,
    \sw_170_module_data_in[5] ,
    \sw_170_module_data_in[4] ,
    \sw_170_module_data_in[3] ,
    \sw_170_module_data_in[2] ,
    \sw_170_module_data_in[1] ,
    \sw_170_module_data_in[0] }),
    .module_data_out({\sw_170_module_data_out[7] ,
    \sw_170_module_data_out[6] ,
    \sw_170_module_data_out[5] ,
    \sw_170_module_data_out[4] ,
    \sw_170_module_data_out[3] ,
    \sw_170_module_data_out[2] ,
    \sw_170_module_data_out[1] ,
    \sw_170_module_data_out[0] }));
 scanchain scanchain_171 (.clk_in(sw_170_clk_out),
    .clk_out(sw_171_clk_out),
    .data_in(sw_170_data_out),
    .data_out(sw_171_data_out),
    .latch_enable_in(sw_170_latch_out),
    .latch_enable_out(sw_171_latch_out),
    .scan_select_in(sw_170_scan_out),
    .scan_select_out(sw_171_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_171_module_data_in[7] ,
    \sw_171_module_data_in[6] ,
    \sw_171_module_data_in[5] ,
    \sw_171_module_data_in[4] ,
    \sw_171_module_data_in[3] ,
    \sw_171_module_data_in[2] ,
    \sw_171_module_data_in[1] ,
    \sw_171_module_data_in[0] }),
    .module_data_out({\sw_171_module_data_out[7] ,
    \sw_171_module_data_out[6] ,
    \sw_171_module_data_out[5] ,
    \sw_171_module_data_out[4] ,
    \sw_171_module_data_out[3] ,
    \sw_171_module_data_out[2] ,
    \sw_171_module_data_out[1] ,
    \sw_171_module_data_out[0] }));
 scanchain scanchain_172 (.clk_in(sw_171_clk_out),
    .clk_out(sw_172_clk_out),
    .data_in(sw_171_data_out),
    .data_out(sw_172_data_out),
    .latch_enable_in(sw_171_latch_out),
    .latch_enable_out(sw_172_latch_out),
    .scan_select_in(sw_171_scan_out),
    .scan_select_out(sw_172_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_172_module_data_in[7] ,
    \sw_172_module_data_in[6] ,
    \sw_172_module_data_in[5] ,
    \sw_172_module_data_in[4] ,
    \sw_172_module_data_in[3] ,
    \sw_172_module_data_in[2] ,
    \sw_172_module_data_in[1] ,
    \sw_172_module_data_in[0] }),
    .module_data_out({\sw_172_module_data_out[7] ,
    \sw_172_module_data_out[6] ,
    \sw_172_module_data_out[5] ,
    \sw_172_module_data_out[4] ,
    \sw_172_module_data_out[3] ,
    \sw_172_module_data_out[2] ,
    \sw_172_module_data_out[1] ,
    \sw_172_module_data_out[0] }));
 scanchain scanchain_173 (.clk_in(sw_172_clk_out),
    .clk_out(sw_173_clk_out),
    .data_in(sw_172_data_out),
    .data_out(sw_173_data_out),
    .latch_enable_in(sw_172_latch_out),
    .latch_enable_out(sw_173_latch_out),
    .scan_select_in(sw_172_scan_out),
    .scan_select_out(sw_173_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_173_module_data_in[7] ,
    \sw_173_module_data_in[6] ,
    \sw_173_module_data_in[5] ,
    \sw_173_module_data_in[4] ,
    \sw_173_module_data_in[3] ,
    \sw_173_module_data_in[2] ,
    \sw_173_module_data_in[1] ,
    \sw_173_module_data_in[0] }),
    .module_data_out({\sw_173_module_data_out[7] ,
    \sw_173_module_data_out[6] ,
    \sw_173_module_data_out[5] ,
    \sw_173_module_data_out[4] ,
    \sw_173_module_data_out[3] ,
    \sw_173_module_data_out[2] ,
    \sw_173_module_data_out[1] ,
    \sw_173_module_data_out[0] }));
 scanchain scanchain_174 (.clk_in(sw_173_clk_out),
    .clk_out(sw_174_clk_out),
    .data_in(sw_173_data_out),
    .data_out(sw_174_data_out),
    .latch_enable_in(sw_173_latch_out),
    .latch_enable_out(sw_174_latch_out),
    .scan_select_in(sw_173_scan_out),
    .scan_select_out(sw_174_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_174_module_data_in[7] ,
    \sw_174_module_data_in[6] ,
    \sw_174_module_data_in[5] ,
    \sw_174_module_data_in[4] ,
    \sw_174_module_data_in[3] ,
    \sw_174_module_data_in[2] ,
    \sw_174_module_data_in[1] ,
    \sw_174_module_data_in[0] }),
    .module_data_out({\sw_174_module_data_out[7] ,
    \sw_174_module_data_out[6] ,
    \sw_174_module_data_out[5] ,
    \sw_174_module_data_out[4] ,
    \sw_174_module_data_out[3] ,
    \sw_174_module_data_out[2] ,
    \sw_174_module_data_out[1] ,
    \sw_174_module_data_out[0] }));
 scanchain scanchain_175 (.clk_in(sw_174_clk_out),
    .clk_out(sw_175_clk_out),
    .data_in(sw_174_data_out),
    .data_out(sw_175_data_out),
    .latch_enable_in(sw_174_latch_out),
    .latch_enable_out(sw_175_latch_out),
    .scan_select_in(sw_174_scan_out),
    .scan_select_out(sw_175_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_175_module_data_in[7] ,
    \sw_175_module_data_in[6] ,
    \sw_175_module_data_in[5] ,
    \sw_175_module_data_in[4] ,
    \sw_175_module_data_in[3] ,
    \sw_175_module_data_in[2] ,
    \sw_175_module_data_in[1] ,
    \sw_175_module_data_in[0] }),
    .module_data_out({\sw_175_module_data_out[7] ,
    \sw_175_module_data_out[6] ,
    \sw_175_module_data_out[5] ,
    \sw_175_module_data_out[4] ,
    \sw_175_module_data_out[3] ,
    \sw_175_module_data_out[2] ,
    \sw_175_module_data_out[1] ,
    \sw_175_module_data_out[0] }));
 scanchain scanchain_176 (.clk_in(sw_175_clk_out),
    .clk_out(sw_176_clk_out),
    .data_in(sw_175_data_out),
    .data_out(sw_176_data_out),
    .latch_enable_in(sw_175_latch_out),
    .latch_enable_out(sw_176_latch_out),
    .scan_select_in(sw_175_scan_out),
    .scan_select_out(sw_176_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_176_module_data_in[7] ,
    \sw_176_module_data_in[6] ,
    \sw_176_module_data_in[5] ,
    \sw_176_module_data_in[4] ,
    \sw_176_module_data_in[3] ,
    \sw_176_module_data_in[2] ,
    \sw_176_module_data_in[1] ,
    \sw_176_module_data_in[0] }),
    .module_data_out({\sw_176_module_data_out[7] ,
    \sw_176_module_data_out[6] ,
    \sw_176_module_data_out[5] ,
    \sw_176_module_data_out[4] ,
    \sw_176_module_data_out[3] ,
    \sw_176_module_data_out[2] ,
    \sw_176_module_data_out[1] ,
    \sw_176_module_data_out[0] }));
 scanchain scanchain_177 (.clk_in(sw_176_clk_out),
    .clk_out(sw_177_clk_out),
    .data_in(sw_176_data_out),
    .data_out(sw_177_data_out),
    .latch_enable_in(sw_176_latch_out),
    .latch_enable_out(sw_177_latch_out),
    .scan_select_in(sw_176_scan_out),
    .scan_select_out(sw_177_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_177_module_data_in[7] ,
    \sw_177_module_data_in[6] ,
    \sw_177_module_data_in[5] ,
    \sw_177_module_data_in[4] ,
    \sw_177_module_data_in[3] ,
    \sw_177_module_data_in[2] ,
    \sw_177_module_data_in[1] ,
    \sw_177_module_data_in[0] }),
    .module_data_out({\sw_177_module_data_out[7] ,
    \sw_177_module_data_out[6] ,
    \sw_177_module_data_out[5] ,
    \sw_177_module_data_out[4] ,
    \sw_177_module_data_out[3] ,
    \sw_177_module_data_out[2] ,
    \sw_177_module_data_out[1] ,
    \sw_177_module_data_out[0] }));
 scanchain scanchain_178 (.clk_in(sw_177_clk_out),
    .clk_out(sw_178_clk_out),
    .data_in(sw_177_data_out),
    .data_out(sw_178_data_out),
    .latch_enable_in(sw_177_latch_out),
    .latch_enable_out(sw_178_latch_out),
    .scan_select_in(sw_177_scan_out),
    .scan_select_out(sw_178_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_178_module_data_in[7] ,
    \sw_178_module_data_in[6] ,
    \sw_178_module_data_in[5] ,
    \sw_178_module_data_in[4] ,
    \sw_178_module_data_in[3] ,
    \sw_178_module_data_in[2] ,
    \sw_178_module_data_in[1] ,
    \sw_178_module_data_in[0] }),
    .module_data_out({\sw_178_module_data_out[7] ,
    \sw_178_module_data_out[6] ,
    \sw_178_module_data_out[5] ,
    \sw_178_module_data_out[4] ,
    \sw_178_module_data_out[3] ,
    \sw_178_module_data_out[2] ,
    \sw_178_module_data_out[1] ,
    \sw_178_module_data_out[0] }));
 scanchain scanchain_179 (.clk_in(sw_178_clk_out),
    .clk_out(sw_179_clk_out),
    .data_in(sw_178_data_out),
    .data_out(sw_179_data_out),
    .latch_enable_in(sw_178_latch_out),
    .latch_enable_out(sw_179_latch_out),
    .scan_select_in(sw_178_scan_out),
    .scan_select_out(sw_179_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_179_module_data_in[7] ,
    \sw_179_module_data_in[6] ,
    \sw_179_module_data_in[5] ,
    \sw_179_module_data_in[4] ,
    \sw_179_module_data_in[3] ,
    \sw_179_module_data_in[2] ,
    \sw_179_module_data_in[1] ,
    \sw_179_module_data_in[0] }),
    .module_data_out({\sw_179_module_data_out[7] ,
    \sw_179_module_data_out[6] ,
    \sw_179_module_data_out[5] ,
    \sw_179_module_data_out[4] ,
    \sw_179_module_data_out[3] ,
    \sw_179_module_data_out[2] ,
    \sw_179_module_data_out[1] ,
    \sw_179_module_data_out[0] }));
 scanchain scanchain_180 (.clk_in(sw_179_clk_out),
    .clk_out(sw_180_clk_out),
    .data_in(sw_179_data_out),
    .data_out(sw_180_data_out),
    .latch_enable_in(sw_179_latch_out),
    .latch_enable_out(sw_180_latch_out),
    .scan_select_in(sw_179_scan_out),
    .scan_select_out(sw_180_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_180_module_data_in[7] ,
    \sw_180_module_data_in[6] ,
    \sw_180_module_data_in[5] ,
    \sw_180_module_data_in[4] ,
    \sw_180_module_data_in[3] ,
    \sw_180_module_data_in[2] ,
    \sw_180_module_data_in[1] ,
    \sw_180_module_data_in[0] }),
    .module_data_out({\sw_180_module_data_out[7] ,
    \sw_180_module_data_out[6] ,
    \sw_180_module_data_out[5] ,
    \sw_180_module_data_out[4] ,
    \sw_180_module_data_out[3] ,
    \sw_180_module_data_out[2] ,
    \sw_180_module_data_out[1] ,
    \sw_180_module_data_out[0] }));
 scanchain scanchain_181 (.clk_in(sw_180_clk_out),
    .clk_out(sw_181_clk_out),
    .data_in(sw_180_data_out),
    .data_out(sw_181_data_out),
    .latch_enable_in(sw_180_latch_out),
    .latch_enable_out(sw_181_latch_out),
    .scan_select_in(sw_180_scan_out),
    .scan_select_out(sw_181_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_181_module_data_in[7] ,
    \sw_181_module_data_in[6] ,
    \sw_181_module_data_in[5] ,
    \sw_181_module_data_in[4] ,
    \sw_181_module_data_in[3] ,
    \sw_181_module_data_in[2] ,
    \sw_181_module_data_in[1] ,
    \sw_181_module_data_in[0] }),
    .module_data_out({\sw_181_module_data_out[7] ,
    \sw_181_module_data_out[6] ,
    \sw_181_module_data_out[5] ,
    \sw_181_module_data_out[4] ,
    \sw_181_module_data_out[3] ,
    \sw_181_module_data_out[2] ,
    \sw_181_module_data_out[1] ,
    \sw_181_module_data_out[0] }));
 scanchain scanchain_182 (.clk_in(sw_181_clk_out),
    .clk_out(sw_182_clk_out),
    .data_in(sw_181_data_out),
    .data_out(sw_182_data_out),
    .latch_enable_in(sw_181_latch_out),
    .latch_enable_out(sw_182_latch_out),
    .scan_select_in(sw_181_scan_out),
    .scan_select_out(sw_182_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_182_module_data_in[7] ,
    \sw_182_module_data_in[6] ,
    \sw_182_module_data_in[5] ,
    \sw_182_module_data_in[4] ,
    \sw_182_module_data_in[3] ,
    \sw_182_module_data_in[2] ,
    \sw_182_module_data_in[1] ,
    \sw_182_module_data_in[0] }),
    .module_data_out({\sw_182_module_data_out[7] ,
    \sw_182_module_data_out[6] ,
    \sw_182_module_data_out[5] ,
    \sw_182_module_data_out[4] ,
    \sw_182_module_data_out[3] ,
    \sw_182_module_data_out[2] ,
    \sw_182_module_data_out[1] ,
    \sw_182_module_data_out[0] }));
 scanchain scanchain_183 (.clk_in(sw_182_clk_out),
    .clk_out(sw_183_clk_out),
    .data_in(sw_182_data_out),
    .data_out(sw_183_data_out),
    .latch_enable_in(sw_182_latch_out),
    .latch_enable_out(sw_183_latch_out),
    .scan_select_in(sw_182_scan_out),
    .scan_select_out(sw_183_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_183_module_data_in[7] ,
    \sw_183_module_data_in[6] ,
    \sw_183_module_data_in[5] ,
    \sw_183_module_data_in[4] ,
    \sw_183_module_data_in[3] ,
    \sw_183_module_data_in[2] ,
    \sw_183_module_data_in[1] ,
    \sw_183_module_data_in[0] }),
    .module_data_out({\sw_183_module_data_out[7] ,
    \sw_183_module_data_out[6] ,
    \sw_183_module_data_out[5] ,
    \sw_183_module_data_out[4] ,
    \sw_183_module_data_out[3] ,
    \sw_183_module_data_out[2] ,
    \sw_183_module_data_out[1] ,
    \sw_183_module_data_out[0] }));
 scanchain scanchain_184 (.clk_in(sw_183_clk_out),
    .clk_out(sw_184_clk_out),
    .data_in(sw_183_data_out),
    .data_out(sw_184_data_out),
    .latch_enable_in(sw_183_latch_out),
    .latch_enable_out(sw_184_latch_out),
    .scan_select_in(sw_183_scan_out),
    .scan_select_out(sw_184_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_184_module_data_in[7] ,
    \sw_184_module_data_in[6] ,
    \sw_184_module_data_in[5] ,
    \sw_184_module_data_in[4] ,
    \sw_184_module_data_in[3] ,
    \sw_184_module_data_in[2] ,
    \sw_184_module_data_in[1] ,
    \sw_184_module_data_in[0] }),
    .module_data_out({\sw_184_module_data_out[7] ,
    \sw_184_module_data_out[6] ,
    \sw_184_module_data_out[5] ,
    \sw_184_module_data_out[4] ,
    \sw_184_module_data_out[3] ,
    \sw_184_module_data_out[2] ,
    \sw_184_module_data_out[1] ,
    \sw_184_module_data_out[0] }));
 scanchain scanchain_185 (.clk_in(sw_184_clk_out),
    .clk_out(sw_185_clk_out),
    .data_in(sw_184_data_out),
    .data_out(sw_185_data_out),
    .latch_enable_in(sw_184_latch_out),
    .latch_enable_out(sw_185_latch_out),
    .scan_select_in(sw_184_scan_out),
    .scan_select_out(sw_185_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_185_module_data_in[7] ,
    \sw_185_module_data_in[6] ,
    \sw_185_module_data_in[5] ,
    \sw_185_module_data_in[4] ,
    \sw_185_module_data_in[3] ,
    \sw_185_module_data_in[2] ,
    \sw_185_module_data_in[1] ,
    \sw_185_module_data_in[0] }),
    .module_data_out({\sw_185_module_data_out[7] ,
    \sw_185_module_data_out[6] ,
    \sw_185_module_data_out[5] ,
    \sw_185_module_data_out[4] ,
    \sw_185_module_data_out[3] ,
    \sw_185_module_data_out[2] ,
    \sw_185_module_data_out[1] ,
    \sw_185_module_data_out[0] }));
 scanchain scanchain_186 (.clk_in(sw_185_clk_out),
    .clk_out(sw_186_clk_out),
    .data_in(sw_185_data_out),
    .data_out(sw_186_data_out),
    .latch_enable_in(sw_185_latch_out),
    .latch_enable_out(sw_186_latch_out),
    .scan_select_in(sw_185_scan_out),
    .scan_select_out(sw_186_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_186_module_data_in[7] ,
    \sw_186_module_data_in[6] ,
    \sw_186_module_data_in[5] ,
    \sw_186_module_data_in[4] ,
    \sw_186_module_data_in[3] ,
    \sw_186_module_data_in[2] ,
    \sw_186_module_data_in[1] ,
    \sw_186_module_data_in[0] }),
    .module_data_out({\sw_186_module_data_out[7] ,
    \sw_186_module_data_out[6] ,
    \sw_186_module_data_out[5] ,
    \sw_186_module_data_out[4] ,
    \sw_186_module_data_out[3] ,
    \sw_186_module_data_out[2] ,
    \sw_186_module_data_out[1] ,
    \sw_186_module_data_out[0] }));
 scanchain scanchain_187 (.clk_in(sw_186_clk_out),
    .clk_out(sw_187_clk_out),
    .data_in(sw_186_data_out),
    .data_out(sw_187_data_out),
    .latch_enable_in(sw_186_latch_out),
    .latch_enable_out(sw_187_latch_out),
    .scan_select_in(sw_186_scan_out),
    .scan_select_out(sw_187_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_187_module_data_in[7] ,
    \sw_187_module_data_in[6] ,
    \sw_187_module_data_in[5] ,
    \sw_187_module_data_in[4] ,
    \sw_187_module_data_in[3] ,
    \sw_187_module_data_in[2] ,
    \sw_187_module_data_in[1] ,
    \sw_187_module_data_in[0] }),
    .module_data_out({\sw_187_module_data_out[7] ,
    \sw_187_module_data_out[6] ,
    \sw_187_module_data_out[5] ,
    \sw_187_module_data_out[4] ,
    \sw_187_module_data_out[3] ,
    \sw_187_module_data_out[2] ,
    \sw_187_module_data_out[1] ,
    \sw_187_module_data_out[0] }));
 scanchain scanchain_188 (.clk_in(sw_187_clk_out),
    .clk_out(sw_188_clk_out),
    .data_in(sw_187_data_out),
    .data_out(sw_188_data_out),
    .latch_enable_in(sw_187_latch_out),
    .latch_enable_out(sw_188_latch_out),
    .scan_select_in(sw_187_scan_out),
    .scan_select_out(sw_188_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_188_module_data_in[7] ,
    \sw_188_module_data_in[6] ,
    \sw_188_module_data_in[5] ,
    \sw_188_module_data_in[4] ,
    \sw_188_module_data_in[3] ,
    \sw_188_module_data_in[2] ,
    \sw_188_module_data_in[1] ,
    \sw_188_module_data_in[0] }),
    .module_data_out({\sw_188_module_data_out[7] ,
    \sw_188_module_data_out[6] ,
    \sw_188_module_data_out[5] ,
    \sw_188_module_data_out[4] ,
    \sw_188_module_data_out[3] ,
    \sw_188_module_data_out[2] ,
    \sw_188_module_data_out[1] ,
    \sw_188_module_data_out[0] }));
 scanchain scanchain_189 (.clk_in(sw_188_clk_out),
    .clk_out(sw_189_clk_out),
    .data_in(sw_188_data_out),
    .data_out(sw_189_data_out),
    .latch_enable_in(sw_188_latch_out),
    .latch_enable_out(sw_189_latch_out),
    .scan_select_in(sw_188_scan_out),
    .scan_select_out(sw_189_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_189_module_data_in[7] ,
    \sw_189_module_data_in[6] ,
    \sw_189_module_data_in[5] ,
    \sw_189_module_data_in[4] ,
    \sw_189_module_data_in[3] ,
    \sw_189_module_data_in[2] ,
    \sw_189_module_data_in[1] ,
    \sw_189_module_data_in[0] }),
    .module_data_out({\sw_189_module_data_out[7] ,
    \sw_189_module_data_out[6] ,
    \sw_189_module_data_out[5] ,
    \sw_189_module_data_out[4] ,
    \sw_189_module_data_out[3] ,
    \sw_189_module_data_out[2] ,
    \sw_189_module_data_out[1] ,
    \sw_189_module_data_out[0] }));
 scanchain scanchain_190 (.clk_in(sw_189_clk_out),
    .clk_out(sw_190_clk_out),
    .data_in(sw_189_data_out),
    .data_out(sw_190_data_out),
    .latch_enable_in(sw_189_latch_out),
    .latch_enable_out(sw_190_latch_out),
    .scan_select_in(sw_189_scan_out),
    .scan_select_out(sw_190_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_190_module_data_in[7] ,
    \sw_190_module_data_in[6] ,
    \sw_190_module_data_in[5] ,
    \sw_190_module_data_in[4] ,
    \sw_190_module_data_in[3] ,
    \sw_190_module_data_in[2] ,
    \sw_190_module_data_in[1] ,
    \sw_190_module_data_in[0] }),
    .module_data_out({\sw_190_module_data_out[7] ,
    \sw_190_module_data_out[6] ,
    \sw_190_module_data_out[5] ,
    \sw_190_module_data_out[4] ,
    \sw_190_module_data_out[3] ,
    \sw_190_module_data_out[2] ,
    \sw_190_module_data_out[1] ,
    \sw_190_module_data_out[0] }));
 scanchain scanchain_191 (.clk_in(sw_190_clk_out),
    .clk_out(sw_191_clk_out),
    .data_in(sw_190_data_out),
    .data_out(sw_191_data_out),
    .latch_enable_in(sw_190_latch_out),
    .latch_enable_out(sw_191_latch_out),
    .scan_select_in(sw_190_scan_out),
    .scan_select_out(sw_191_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_191_module_data_in[7] ,
    \sw_191_module_data_in[6] ,
    \sw_191_module_data_in[5] ,
    \sw_191_module_data_in[4] ,
    \sw_191_module_data_in[3] ,
    \sw_191_module_data_in[2] ,
    \sw_191_module_data_in[1] ,
    \sw_191_module_data_in[0] }),
    .module_data_out({\sw_191_module_data_out[7] ,
    \sw_191_module_data_out[6] ,
    \sw_191_module_data_out[5] ,
    \sw_191_module_data_out[4] ,
    \sw_191_module_data_out[3] ,
    \sw_191_module_data_out[2] ,
    \sw_191_module_data_out[1] ,
    \sw_191_module_data_out[0] }));
 scanchain scanchain_192 (.clk_in(sw_191_clk_out),
    .clk_out(sw_192_clk_out),
    .data_in(sw_191_data_out),
    .data_out(sw_192_data_out),
    .latch_enable_in(sw_191_latch_out),
    .latch_enable_out(sw_192_latch_out),
    .scan_select_in(sw_191_scan_out),
    .scan_select_out(sw_192_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_192_module_data_in[7] ,
    \sw_192_module_data_in[6] ,
    \sw_192_module_data_in[5] ,
    \sw_192_module_data_in[4] ,
    \sw_192_module_data_in[3] ,
    \sw_192_module_data_in[2] ,
    \sw_192_module_data_in[1] ,
    \sw_192_module_data_in[0] }),
    .module_data_out({\sw_192_module_data_out[7] ,
    \sw_192_module_data_out[6] ,
    \sw_192_module_data_out[5] ,
    \sw_192_module_data_out[4] ,
    \sw_192_module_data_out[3] ,
    \sw_192_module_data_out[2] ,
    \sw_192_module_data_out[1] ,
    \sw_192_module_data_out[0] }));
 scanchain scanchain_193 (.clk_in(sw_192_clk_out),
    .clk_out(sw_193_clk_out),
    .data_in(sw_192_data_out),
    .data_out(sw_193_data_out),
    .latch_enable_in(sw_192_latch_out),
    .latch_enable_out(sw_193_latch_out),
    .scan_select_in(sw_192_scan_out),
    .scan_select_out(sw_193_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_193_module_data_in[7] ,
    \sw_193_module_data_in[6] ,
    \sw_193_module_data_in[5] ,
    \sw_193_module_data_in[4] ,
    \sw_193_module_data_in[3] ,
    \sw_193_module_data_in[2] ,
    \sw_193_module_data_in[1] ,
    \sw_193_module_data_in[0] }),
    .module_data_out({\sw_193_module_data_out[7] ,
    \sw_193_module_data_out[6] ,
    \sw_193_module_data_out[5] ,
    \sw_193_module_data_out[4] ,
    \sw_193_module_data_out[3] ,
    \sw_193_module_data_out[2] ,
    \sw_193_module_data_out[1] ,
    \sw_193_module_data_out[0] }));
 scanchain scanchain_194 (.clk_in(sw_193_clk_out),
    .clk_out(sw_194_clk_out),
    .data_in(sw_193_data_out),
    .data_out(sw_194_data_out),
    .latch_enable_in(sw_193_latch_out),
    .latch_enable_out(sw_194_latch_out),
    .scan_select_in(sw_193_scan_out),
    .scan_select_out(sw_194_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_194_module_data_in[7] ,
    \sw_194_module_data_in[6] ,
    \sw_194_module_data_in[5] ,
    \sw_194_module_data_in[4] ,
    \sw_194_module_data_in[3] ,
    \sw_194_module_data_in[2] ,
    \sw_194_module_data_in[1] ,
    \sw_194_module_data_in[0] }),
    .module_data_out({\sw_194_module_data_out[7] ,
    \sw_194_module_data_out[6] ,
    \sw_194_module_data_out[5] ,
    \sw_194_module_data_out[4] ,
    \sw_194_module_data_out[3] ,
    \sw_194_module_data_out[2] ,
    \sw_194_module_data_out[1] ,
    \sw_194_module_data_out[0] }));
 scanchain scanchain_195 (.clk_in(sw_194_clk_out),
    .clk_out(sw_195_clk_out),
    .data_in(sw_194_data_out),
    .data_out(sw_195_data_out),
    .latch_enable_in(sw_194_latch_out),
    .latch_enable_out(sw_195_latch_out),
    .scan_select_in(sw_194_scan_out),
    .scan_select_out(sw_195_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_195_module_data_in[7] ,
    \sw_195_module_data_in[6] ,
    \sw_195_module_data_in[5] ,
    \sw_195_module_data_in[4] ,
    \sw_195_module_data_in[3] ,
    \sw_195_module_data_in[2] ,
    \sw_195_module_data_in[1] ,
    \sw_195_module_data_in[0] }),
    .module_data_out({\sw_195_module_data_out[7] ,
    \sw_195_module_data_out[6] ,
    \sw_195_module_data_out[5] ,
    \sw_195_module_data_out[4] ,
    \sw_195_module_data_out[3] ,
    \sw_195_module_data_out[2] ,
    \sw_195_module_data_out[1] ,
    \sw_195_module_data_out[0] }));
 scanchain scanchain_196 (.clk_in(sw_195_clk_out),
    .clk_out(sw_196_clk_out),
    .data_in(sw_195_data_out),
    .data_out(sw_196_data_out),
    .latch_enable_in(sw_195_latch_out),
    .latch_enable_out(sw_196_latch_out),
    .scan_select_in(sw_195_scan_out),
    .scan_select_out(sw_196_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_196_module_data_in[7] ,
    \sw_196_module_data_in[6] ,
    \sw_196_module_data_in[5] ,
    \sw_196_module_data_in[4] ,
    \sw_196_module_data_in[3] ,
    \sw_196_module_data_in[2] ,
    \sw_196_module_data_in[1] ,
    \sw_196_module_data_in[0] }),
    .module_data_out({\sw_196_module_data_out[7] ,
    \sw_196_module_data_out[6] ,
    \sw_196_module_data_out[5] ,
    \sw_196_module_data_out[4] ,
    \sw_196_module_data_out[3] ,
    \sw_196_module_data_out[2] ,
    \sw_196_module_data_out[1] ,
    \sw_196_module_data_out[0] }));
 scanchain scanchain_197 (.clk_in(sw_196_clk_out),
    .clk_out(sw_197_clk_out),
    .data_in(sw_196_data_out),
    .data_out(sw_197_data_out),
    .latch_enable_in(sw_196_latch_out),
    .latch_enable_out(sw_197_latch_out),
    .scan_select_in(sw_196_scan_out),
    .scan_select_out(sw_197_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_197_module_data_in[7] ,
    \sw_197_module_data_in[6] ,
    \sw_197_module_data_in[5] ,
    \sw_197_module_data_in[4] ,
    \sw_197_module_data_in[3] ,
    \sw_197_module_data_in[2] ,
    \sw_197_module_data_in[1] ,
    \sw_197_module_data_in[0] }),
    .module_data_out({\sw_197_module_data_out[7] ,
    \sw_197_module_data_out[6] ,
    \sw_197_module_data_out[5] ,
    \sw_197_module_data_out[4] ,
    \sw_197_module_data_out[3] ,
    \sw_197_module_data_out[2] ,
    \sw_197_module_data_out[1] ,
    \sw_197_module_data_out[0] }));
 scanchain scanchain_198 (.clk_in(sw_197_clk_out),
    .clk_out(sw_198_clk_out),
    .data_in(sw_197_data_out),
    .data_out(sw_198_data_out),
    .latch_enable_in(sw_197_latch_out),
    .latch_enable_out(sw_198_latch_out),
    .scan_select_in(sw_197_scan_out),
    .scan_select_out(sw_198_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_198_module_data_in[7] ,
    \sw_198_module_data_in[6] ,
    \sw_198_module_data_in[5] ,
    \sw_198_module_data_in[4] ,
    \sw_198_module_data_in[3] ,
    \sw_198_module_data_in[2] ,
    \sw_198_module_data_in[1] ,
    \sw_198_module_data_in[0] }),
    .module_data_out({\sw_198_module_data_out[7] ,
    \sw_198_module_data_out[6] ,
    \sw_198_module_data_out[5] ,
    \sw_198_module_data_out[4] ,
    \sw_198_module_data_out[3] ,
    \sw_198_module_data_out[2] ,
    \sw_198_module_data_out[1] ,
    \sw_198_module_data_out[0] }));
 scanchain scanchain_199 (.clk_in(sw_198_clk_out),
    .clk_out(sw_199_clk_out),
    .data_in(sw_198_data_out),
    .data_out(sw_199_data_out),
    .latch_enable_in(sw_198_latch_out),
    .latch_enable_out(sw_199_latch_out),
    .scan_select_in(sw_198_scan_out),
    .scan_select_out(sw_199_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_199_module_data_in[7] ,
    \sw_199_module_data_in[6] ,
    \sw_199_module_data_in[5] ,
    \sw_199_module_data_in[4] ,
    \sw_199_module_data_in[3] ,
    \sw_199_module_data_in[2] ,
    \sw_199_module_data_in[1] ,
    \sw_199_module_data_in[0] }),
    .module_data_out({\sw_199_module_data_out[7] ,
    \sw_199_module_data_out[6] ,
    \sw_199_module_data_out[5] ,
    \sw_199_module_data_out[4] ,
    \sw_199_module_data_out[3] ,
    \sw_199_module_data_out[2] ,
    \sw_199_module_data_out[1] ,
    \sw_199_module_data_out[0] }));
 scanchain scanchain_200 (.clk_in(sw_199_clk_out),
    .clk_out(sw_200_clk_out),
    .data_in(sw_199_data_out),
    .data_out(sw_200_data_out),
    .latch_enable_in(sw_199_latch_out),
    .latch_enable_out(sw_200_latch_out),
    .scan_select_in(sw_199_scan_out),
    .scan_select_out(sw_200_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_200_module_data_in[7] ,
    \sw_200_module_data_in[6] ,
    \sw_200_module_data_in[5] ,
    \sw_200_module_data_in[4] ,
    \sw_200_module_data_in[3] ,
    \sw_200_module_data_in[2] ,
    \sw_200_module_data_in[1] ,
    \sw_200_module_data_in[0] }),
    .module_data_out({\sw_200_module_data_out[7] ,
    \sw_200_module_data_out[6] ,
    \sw_200_module_data_out[5] ,
    \sw_200_module_data_out[4] ,
    \sw_200_module_data_out[3] ,
    \sw_200_module_data_out[2] ,
    \sw_200_module_data_out[1] ,
    \sw_200_module_data_out[0] }));
 scanchain scanchain_201 (.clk_in(sw_200_clk_out),
    .clk_out(sw_201_clk_out),
    .data_in(sw_200_data_out),
    .data_out(sw_201_data_out),
    .latch_enable_in(sw_200_latch_out),
    .latch_enable_out(sw_201_latch_out),
    .scan_select_in(sw_200_scan_out),
    .scan_select_out(sw_201_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_201_module_data_in[7] ,
    \sw_201_module_data_in[6] ,
    \sw_201_module_data_in[5] ,
    \sw_201_module_data_in[4] ,
    \sw_201_module_data_in[3] ,
    \sw_201_module_data_in[2] ,
    \sw_201_module_data_in[1] ,
    \sw_201_module_data_in[0] }),
    .module_data_out({\sw_201_module_data_out[7] ,
    \sw_201_module_data_out[6] ,
    \sw_201_module_data_out[5] ,
    \sw_201_module_data_out[4] ,
    \sw_201_module_data_out[3] ,
    \sw_201_module_data_out[2] ,
    \sw_201_module_data_out[1] ,
    \sw_201_module_data_out[0] }));
 scanchain scanchain_202 (.clk_in(sw_201_clk_out),
    .clk_out(sw_202_clk_out),
    .data_in(sw_201_data_out),
    .data_out(sw_202_data_out),
    .latch_enable_in(sw_201_latch_out),
    .latch_enable_out(sw_202_latch_out),
    .scan_select_in(sw_201_scan_out),
    .scan_select_out(sw_202_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_202_module_data_in[7] ,
    \sw_202_module_data_in[6] ,
    \sw_202_module_data_in[5] ,
    \sw_202_module_data_in[4] ,
    \sw_202_module_data_in[3] ,
    \sw_202_module_data_in[2] ,
    \sw_202_module_data_in[1] ,
    \sw_202_module_data_in[0] }),
    .module_data_out({\sw_202_module_data_out[7] ,
    \sw_202_module_data_out[6] ,
    \sw_202_module_data_out[5] ,
    \sw_202_module_data_out[4] ,
    \sw_202_module_data_out[3] ,
    \sw_202_module_data_out[2] ,
    \sw_202_module_data_out[1] ,
    \sw_202_module_data_out[0] }));
 scanchain scanchain_203 (.clk_in(sw_202_clk_out),
    .clk_out(sw_203_clk_out),
    .data_in(sw_202_data_out),
    .data_out(sw_203_data_out),
    .latch_enable_in(sw_202_latch_out),
    .latch_enable_out(sw_203_latch_out),
    .scan_select_in(sw_202_scan_out),
    .scan_select_out(sw_203_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_203_module_data_in[7] ,
    \sw_203_module_data_in[6] ,
    \sw_203_module_data_in[5] ,
    \sw_203_module_data_in[4] ,
    \sw_203_module_data_in[3] ,
    \sw_203_module_data_in[2] ,
    \sw_203_module_data_in[1] ,
    \sw_203_module_data_in[0] }),
    .module_data_out({\sw_203_module_data_out[7] ,
    \sw_203_module_data_out[6] ,
    \sw_203_module_data_out[5] ,
    \sw_203_module_data_out[4] ,
    \sw_203_module_data_out[3] ,
    \sw_203_module_data_out[2] ,
    \sw_203_module_data_out[1] ,
    \sw_203_module_data_out[0] }));
 scanchain scanchain_204 (.clk_in(sw_203_clk_out),
    .clk_out(sw_204_clk_out),
    .data_in(sw_203_data_out),
    .data_out(sw_204_data_out),
    .latch_enable_in(sw_203_latch_out),
    .latch_enable_out(sw_204_latch_out),
    .scan_select_in(sw_203_scan_out),
    .scan_select_out(sw_204_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_204_module_data_in[7] ,
    \sw_204_module_data_in[6] ,
    \sw_204_module_data_in[5] ,
    \sw_204_module_data_in[4] ,
    \sw_204_module_data_in[3] ,
    \sw_204_module_data_in[2] ,
    \sw_204_module_data_in[1] ,
    \sw_204_module_data_in[0] }),
    .module_data_out({\sw_204_module_data_out[7] ,
    \sw_204_module_data_out[6] ,
    \sw_204_module_data_out[5] ,
    \sw_204_module_data_out[4] ,
    \sw_204_module_data_out[3] ,
    \sw_204_module_data_out[2] ,
    \sw_204_module_data_out[1] ,
    \sw_204_module_data_out[0] }));
 scanchain scanchain_205 (.clk_in(sw_204_clk_out),
    .clk_out(sw_205_clk_out),
    .data_in(sw_204_data_out),
    .data_out(sw_205_data_out),
    .latch_enable_in(sw_204_latch_out),
    .latch_enable_out(sw_205_latch_out),
    .scan_select_in(sw_204_scan_out),
    .scan_select_out(sw_205_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_205_module_data_in[7] ,
    \sw_205_module_data_in[6] ,
    \sw_205_module_data_in[5] ,
    \sw_205_module_data_in[4] ,
    \sw_205_module_data_in[3] ,
    \sw_205_module_data_in[2] ,
    \sw_205_module_data_in[1] ,
    \sw_205_module_data_in[0] }),
    .module_data_out({\sw_205_module_data_out[7] ,
    \sw_205_module_data_out[6] ,
    \sw_205_module_data_out[5] ,
    \sw_205_module_data_out[4] ,
    \sw_205_module_data_out[3] ,
    \sw_205_module_data_out[2] ,
    \sw_205_module_data_out[1] ,
    \sw_205_module_data_out[0] }));
 scanchain scanchain_206 (.clk_in(sw_205_clk_out),
    .clk_out(sw_206_clk_out),
    .data_in(sw_205_data_out),
    .data_out(sw_206_data_out),
    .latch_enable_in(sw_205_latch_out),
    .latch_enable_out(sw_206_latch_out),
    .scan_select_in(sw_205_scan_out),
    .scan_select_out(sw_206_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_206_module_data_in[7] ,
    \sw_206_module_data_in[6] ,
    \sw_206_module_data_in[5] ,
    \sw_206_module_data_in[4] ,
    \sw_206_module_data_in[3] ,
    \sw_206_module_data_in[2] ,
    \sw_206_module_data_in[1] ,
    \sw_206_module_data_in[0] }),
    .module_data_out({\sw_206_module_data_out[7] ,
    \sw_206_module_data_out[6] ,
    \sw_206_module_data_out[5] ,
    \sw_206_module_data_out[4] ,
    \sw_206_module_data_out[3] ,
    \sw_206_module_data_out[2] ,
    \sw_206_module_data_out[1] ,
    \sw_206_module_data_out[0] }));
 scanchain scanchain_207 (.clk_in(sw_206_clk_out),
    .clk_out(sw_207_clk_out),
    .data_in(sw_206_data_out),
    .data_out(sw_207_data_out),
    .latch_enable_in(sw_206_latch_out),
    .latch_enable_out(sw_207_latch_out),
    .scan_select_in(sw_206_scan_out),
    .scan_select_out(sw_207_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_207_module_data_in[7] ,
    \sw_207_module_data_in[6] ,
    \sw_207_module_data_in[5] ,
    \sw_207_module_data_in[4] ,
    \sw_207_module_data_in[3] ,
    \sw_207_module_data_in[2] ,
    \sw_207_module_data_in[1] ,
    \sw_207_module_data_in[0] }),
    .module_data_out({\sw_207_module_data_out[7] ,
    \sw_207_module_data_out[6] ,
    \sw_207_module_data_out[5] ,
    \sw_207_module_data_out[4] ,
    \sw_207_module_data_out[3] ,
    \sw_207_module_data_out[2] ,
    \sw_207_module_data_out[1] ,
    \sw_207_module_data_out[0] }));
 scanchain scanchain_208 (.clk_in(sw_207_clk_out),
    .clk_out(sw_208_clk_out),
    .data_in(sw_207_data_out),
    .data_out(sw_208_data_out),
    .latch_enable_in(sw_207_latch_out),
    .latch_enable_out(sw_208_latch_out),
    .scan_select_in(sw_207_scan_out),
    .scan_select_out(sw_208_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_208_module_data_in[7] ,
    \sw_208_module_data_in[6] ,
    \sw_208_module_data_in[5] ,
    \sw_208_module_data_in[4] ,
    \sw_208_module_data_in[3] ,
    \sw_208_module_data_in[2] ,
    \sw_208_module_data_in[1] ,
    \sw_208_module_data_in[0] }),
    .module_data_out({\sw_208_module_data_out[7] ,
    \sw_208_module_data_out[6] ,
    \sw_208_module_data_out[5] ,
    \sw_208_module_data_out[4] ,
    \sw_208_module_data_out[3] ,
    \sw_208_module_data_out[2] ,
    \sw_208_module_data_out[1] ,
    \sw_208_module_data_out[0] }));
 scanchain scanchain_209 (.clk_in(sw_208_clk_out),
    .clk_out(sw_209_clk_out),
    .data_in(sw_208_data_out),
    .data_out(sw_209_data_out),
    .latch_enable_in(sw_208_latch_out),
    .latch_enable_out(sw_209_latch_out),
    .scan_select_in(sw_208_scan_out),
    .scan_select_out(sw_209_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_209_module_data_in[7] ,
    \sw_209_module_data_in[6] ,
    \sw_209_module_data_in[5] ,
    \sw_209_module_data_in[4] ,
    \sw_209_module_data_in[3] ,
    \sw_209_module_data_in[2] ,
    \sw_209_module_data_in[1] ,
    \sw_209_module_data_in[0] }),
    .module_data_out({\sw_209_module_data_out[7] ,
    \sw_209_module_data_out[6] ,
    \sw_209_module_data_out[5] ,
    \sw_209_module_data_out[4] ,
    \sw_209_module_data_out[3] ,
    \sw_209_module_data_out[2] ,
    \sw_209_module_data_out[1] ,
    \sw_209_module_data_out[0] }));
 scanchain scanchain_210 (.clk_in(sw_209_clk_out),
    .clk_out(sw_210_clk_out),
    .data_in(sw_209_data_out),
    .data_out(sw_210_data_out),
    .latch_enable_in(sw_209_latch_out),
    .latch_enable_out(sw_210_latch_out),
    .scan_select_in(sw_209_scan_out),
    .scan_select_out(sw_210_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_210_module_data_in[7] ,
    \sw_210_module_data_in[6] ,
    \sw_210_module_data_in[5] ,
    \sw_210_module_data_in[4] ,
    \sw_210_module_data_in[3] ,
    \sw_210_module_data_in[2] ,
    \sw_210_module_data_in[1] ,
    \sw_210_module_data_in[0] }),
    .module_data_out({\sw_210_module_data_out[7] ,
    \sw_210_module_data_out[6] ,
    \sw_210_module_data_out[5] ,
    \sw_210_module_data_out[4] ,
    \sw_210_module_data_out[3] ,
    \sw_210_module_data_out[2] ,
    \sw_210_module_data_out[1] ,
    \sw_210_module_data_out[0] }));
 scanchain scanchain_211 (.clk_in(sw_210_clk_out),
    .clk_out(sw_211_clk_out),
    .data_in(sw_210_data_out),
    .data_out(sw_211_data_out),
    .latch_enable_in(sw_210_latch_out),
    .latch_enable_out(sw_211_latch_out),
    .scan_select_in(sw_210_scan_out),
    .scan_select_out(sw_211_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_211_module_data_in[7] ,
    \sw_211_module_data_in[6] ,
    \sw_211_module_data_in[5] ,
    \sw_211_module_data_in[4] ,
    \sw_211_module_data_in[3] ,
    \sw_211_module_data_in[2] ,
    \sw_211_module_data_in[1] ,
    \sw_211_module_data_in[0] }),
    .module_data_out({\sw_211_module_data_out[7] ,
    \sw_211_module_data_out[6] ,
    \sw_211_module_data_out[5] ,
    \sw_211_module_data_out[4] ,
    \sw_211_module_data_out[3] ,
    \sw_211_module_data_out[2] ,
    \sw_211_module_data_out[1] ,
    \sw_211_module_data_out[0] }));
 scanchain scanchain_212 (.clk_in(sw_211_clk_out),
    .clk_out(sw_212_clk_out),
    .data_in(sw_211_data_out),
    .data_out(sw_212_data_out),
    .latch_enable_in(sw_211_latch_out),
    .latch_enable_out(sw_212_latch_out),
    .scan_select_in(sw_211_scan_out),
    .scan_select_out(sw_212_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_212_module_data_in[7] ,
    \sw_212_module_data_in[6] ,
    \sw_212_module_data_in[5] ,
    \sw_212_module_data_in[4] ,
    \sw_212_module_data_in[3] ,
    \sw_212_module_data_in[2] ,
    \sw_212_module_data_in[1] ,
    \sw_212_module_data_in[0] }),
    .module_data_out({\sw_212_module_data_out[7] ,
    \sw_212_module_data_out[6] ,
    \sw_212_module_data_out[5] ,
    \sw_212_module_data_out[4] ,
    \sw_212_module_data_out[3] ,
    \sw_212_module_data_out[2] ,
    \sw_212_module_data_out[1] ,
    \sw_212_module_data_out[0] }));
 scanchain scanchain_213 (.clk_in(sw_212_clk_out),
    .clk_out(sw_213_clk_out),
    .data_in(sw_212_data_out),
    .data_out(sw_213_data_out),
    .latch_enable_in(sw_212_latch_out),
    .latch_enable_out(sw_213_latch_out),
    .scan_select_in(sw_212_scan_out),
    .scan_select_out(sw_213_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_213_module_data_in[7] ,
    \sw_213_module_data_in[6] ,
    \sw_213_module_data_in[5] ,
    \sw_213_module_data_in[4] ,
    \sw_213_module_data_in[3] ,
    \sw_213_module_data_in[2] ,
    \sw_213_module_data_in[1] ,
    \sw_213_module_data_in[0] }),
    .module_data_out({\sw_213_module_data_out[7] ,
    \sw_213_module_data_out[6] ,
    \sw_213_module_data_out[5] ,
    \sw_213_module_data_out[4] ,
    \sw_213_module_data_out[3] ,
    \sw_213_module_data_out[2] ,
    \sw_213_module_data_out[1] ,
    \sw_213_module_data_out[0] }));
 scanchain scanchain_214 (.clk_in(sw_213_clk_out),
    .clk_out(sw_214_clk_out),
    .data_in(sw_213_data_out),
    .data_out(sw_214_data_out),
    .latch_enable_in(sw_213_latch_out),
    .latch_enable_out(sw_214_latch_out),
    .scan_select_in(sw_213_scan_out),
    .scan_select_out(sw_214_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_214_module_data_in[7] ,
    \sw_214_module_data_in[6] ,
    \sw_214_module_data_in[5] ,
    \sw_214_module_data_in[4] ,
    \sw_214_module_data_in[3] ,
    \sw_214_module_data_in[2] ,
    \sw_214_module_data_in[1] ,
    \sw_214_module_data_in[0] }),
    .module_data_out({\sw_214_module_data_out[7] ,
    \sw_214_module_data_out[6] ,
    \sw_214_module_data_out[5] ,
    \sw_214_module_data_out[4] ,
    \sw_214_module_data_out[3] ,
    \sw_214_module_data_out[2] ,
    \sw_214_module_data_out[1] ,
    \sw_214_module_data_out[0] }));
 scanchain scanchain_215 (.clk_in(sw_214_clk_out),
    .clk_out(sw_215_clk_out),
    .data_in(sw_214_data_out),
    .data_out(sw_215_data_out),
    .latch_enable_in(sw_214_latch_out),
    .latch_enable_out(sw_215_latch_out),
    .scan_select_in(sw_214_scan_out),
    .scan_select_out(sw_215_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_215_module_data_in[7] ,
    \sw_215_module_data_in[6] ,
    \sw_215_module_data_in[5] ,
    \sw_215_module_data_in[4] ,
    \sw_215_module_data_in[3] ,
    \sw_215_module_data_in[2] ,
    \sw_215_module_data_in[1] ,
    \sw_215_module_data_in[0] }),
    .module_data_out({\sw_215_module_data_out[7] ,
    \sw_215_module_data_out[6] ,
    \sw_215_module_data_out[5] ,
    \sw_215_module_data_out[4] ,
    \sw_215_module_data_out[3] ,
    \sw_215_module_data_out[2] ,
    \sw_215_module_data_out[1] ,
    \sw_215_module_data_out[0] }));
 scanchain scanchain_216 (.clk_in(sw_215_clk_out),
    .clk_out(sw_216_clk_out),
    .data_in(sw_215_data_out),
    .data_out(sw_216_data_out),
    .latch_enable_in(sw_215_latch_out),
    .latch_enable_out(sw_216_latch_out),
    .scan_select_in(sw_215_scan_out),
    .scan_select_out(sw_216_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_216_module_data_in[7] ,
    \sw_216_module_data_in[6] ,
    \sw_216_module_data_in[5] ,
    \sw_216_module_data_in[4] ,
    \sw_216_module_data_in[3] ,
    \sw_216_module_data_in[2] ,
    \sw_216_module_data_in[1] ,
    \sw_216_module_data_in[0] }),
    .module_data_out({\sw_216_module_data_out[7] ,
    \sw_216_module_data_out[6] ,
    \sw_216_module_data_out[5] ,
    \sw_216_module_data_out[4] ,
    \sw_216_module_data_out[3] ,
    \sw_216_module_data_out[2] ,
    \sw_216_module_data_out[1] ,
    \sw_216_module_data_out[0] }));
 scanchain scanchain_217 (.clk_in(sw_216_clk_out),
    .clk_out(sw_217_clk_out),
    .data_in(sw_216_data_out),
    .data_out(sw_217_data_out),
    .latch_enable_in(sw_216_latch_out),
    .latch_enable_out(sw_217_latch_out),
    .scan_select_in(sw_216_scan_out),
    .scan_select_out(sw_217_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_217_module_data_in[7] ,
    \sw_217_module_data_in[6] ,
    \sw_217_module_data_in[5] ,
    \sw_217_module_data_in[4] ,
    \sw_217_module_data_in[3] ,
    \sw_217_module_data_in[2] ,
    \sw_217_module_data_in[1] ,
    \sw_217_module_data_in[0] }),
    .module_data_out({\sw_217_module_data_out[7] ,
    \sw_217_module_data_out[6] ,
    \sw_217_module_data_out[5] ,
    \sw_217_module_data_out[4] ,
    \sw_217_module_data_out[3] ,
    \sw_217_module_data_out[2] ,
    \sw_217_module_data_out[1] ,
    \sw_217_module_data_out[0] }));
 scanchain scanchain_218 (.clk_in(sw_217_clk_out),
    .clk_out(sw_218_clk_out),
    .data_in(sw_217_data_out),
    .data_out(sw_218_data_out),
    .latch_enable_in(sw_217_latch_out),
    .latch_enable_out(sw_218_latch_out),
    .scan_select_in(sw_217_scan_out),
    .scan_select_out(sw_218_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_218_module_data_in[7] ,
    \sw_218_module_data_in[6] ,
    \sw_218_module_data_in[5] ,
    \sw_218_module_data_in[4] ,
    \sw_218_module_data_in[3] ,
    \sw_218_module_data_in[2] ,
    \sw_218_module_data_in[1] ,
    \sw_218_module_data_in[0] }),
    .module_data_out({\sw_218_module_data_out[7] ,
    \sw_218_module_data_out[6] ,
    \sw_218_module_data_out[5] ,
    \sw_218_module_data_out[4] ,
    \sw_218_module_data_out[3] ,
    \sw_218_module_data_out[2] ,
    \sw_218_module_data_out[1] ,
    \sw_218_module_data_out[0] }));
 scanchain scanchain_219 (.clk_in(sw_218_clk_out),
    .clk_out(sw_219_clk_out),
    .data_in(sw_218_data_out),
    .data_out(sw_219_data_out),
    .latch_enable_in(sw_218_latch_out),
    .latch_enable_out(sw_219_latch_out),
    .scan_select_in(sw_218_scan_out),
    .scan_select_out(sw_219_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_219_module_data_in[7] ,
    \sw_219_module_data_in[6] ,
    \sw_219_module_data_in[5] ,
    \sw_219_module_data_in[4] ,
    \sw_219_module_data_in[3] ,
    \sw_219_module_data_in[2] ,
    \sw_219_module_data_in[1] ,
    \sw_219_module_data_in[0] }),
    .module_data_out({\sw_219_module_data_out[7] ,
    \sw_219_module_data_out[6] ,
    \sw_219_module_data_out[5] ,
    \sw_219_module_data_out[4] ,
    \sw_219_module_data_out[3] ,
    \sw_219_module_data_out[2] ,
    \sw_219_module_data_out[1] ,
    \sw_219_module_data_out[0] }));
 scanchain scanchain_220 (.clk_in(sw_219_clk_out),
    .clk_out(sw_220_clk_out),
    .data_in(sw_219_data_out),
    .data_out(sw_220_data_out),
    .latch_enable_in(sw_219_latch_out),
    .latch_enable_out(sw_220_latch_out),
    .scan_select_in(sw_219_scan_out),
    .scan_select_out(sw_220_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_220_module_data_in[7] ,
    \sw_220_module_data_in[6] ,
    \sw_220_module_data_in[5] ,
    \sw_220_module_data_in[4] ,
    \sw_220_module_data_in[3] ,
    \sw_220_module_data_in[2] ,
    \sw_220_module_data_in[1] ,
    \sw_220_module_data_in[0] }),
    .module_data_out({\sw_220_module_data_out[7] ,
    \sw_220_module_data_out[6] ,
    \sw_220_module_data_out[5] ,
    \sw_220_module_data_out[4] ,
    \sw_220_module_data_out[3] ,
    \sw_220_module_data_out[2] ,
    \sw_220_module_data_out[1] ,
    \sw_220_module_data_out[0] }));
 scanchain scanchain_221 (.clk_in(sw_220_clk_out),
    .clk_out(sw_221_clk_out),
    .data_in(sw_220_data_out),
    .data_out(sw_221_data_out),
    .latch_enable_in(sw_220_latch_out),
    .latch_enable_out(sw_221_latch_out),
    .scan_select_in(sw_220_scan_out),
    .scan_select_out(sw_221_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_221_module_data_in[7] ,
    \sw_221_module_data_in[6] ,
    \sw_221_module_data_in[5] ,
    \sw_221_module_data_in[4] ,
    \sw_221_module_data_in[3] ,
    \sw_221_module_data_in[2] ,
    \sw_221_module_data_in[1] ,
    \sw_221_module_data_in[0] }),
    .module_data_out({\sw_221_module_data_out[7] ,
    \sw_221_module_data_out[6] ,
    \sw_221_module_data_out[5] ,
    \sw_221_module_data_out[4] ,
    \sw_221_module_data_out[3] ,
    \sw_221_module_data_out[2] ,
    \sw_221_module_data_out[1] ,
    \sw_221_module_data_out[0] }));
 scanchain scanchain_222 (.clk_in(sw_221_clk_out),
    .clk_out(sw_222_clk_out),
    .data_in(sw_221_data_out),
    .data_out(sw_222_data_out),
    .latch_enable_in(sw_221_latch_out),
    .latch_enable_out(sw_222_latch_out),
    .scan_select_in(sw_221_scan_out),
    .scan_select_out(sw_222_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_222_module_data_in[7] ,
    \sw_222_module_data_in[6] ,
    \sw_222_module_data_in[5] ,
    \sw_222_module_data_in[4] ,
    \sw_222_module_data_in[3] ,
    \sw_222_module_data_in[2] ,
    \sw_222_module_data_in[1] ,
    \sw_222_module_data_in[0] }),
    .module_data_out({\sw_222_module_data_out[7] ,
    \sw_222_module_data_out[6] ,
    \sw_222_module_data_out[5] ,
    \sw_222_module_data_out[4] ,
    \sw_222_module_data_out[3] ,
    \sw_222_module_data_out[2] ,
    \sw_222_module_data_out[1] ,
    \sw_222_module_data_out[0] }));
 scanchain scanchain_223 (.clk_in(sw_222_clk_out),
    .clk_out(sw_223_clk_out),
    .data_in(sw_222_data_out),
    .data_out(sw_223_data_out),
    .latch_enable_in(sw_222_latch_out),
    .latch_enable_out(sw_223_latch_out),
    .scan_select_in(sw_222_scan_out),
    .scan_select_out(sw_223_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_223_module_data_in[7] ,
    \sw_223_module_data_in[6] ,
    \sw_223_module_data_in[5] ,
    \sw_223_module_data_in[4] ,
    \sw_223_module_data_in[3] ,
    \sw_223_module_data_in[2] ,
    \sw_223_module_data_in[1] ,
    \sw_223_module_data_in[0] }),
    .module_data_out({\sw_223_module_data_out[7] ,
    \sw_223_module_data_out[6] ,
    \sw_223_module_data_out[5] ,
    \sw_223_module_data_out[4] ,
    \sw_223_module_data_out[3] ,
    \sw_223_module_data_out[2] ,
    \sw_223_module_data_out[1] ,
    \sw_223_module_data_out[0] }));
 scanchain scanchain_224 (.clk_in(sw_223_clk_out),
    .clk_out(sw_224_clk_out),
    .data_in(sw_223_data_out),
    .data_out(sw_224_data_out),
    .latch_enable_in(sw_223_latch_out),
    .latch_enable_out(sw_224_latch_out),
    .scan_select_in(sw_223_scan_out),
    .scan_select_out(sw_224_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_224_module_data_in[7] ,
    \sw_224_module_data_in[6] ,
    \sw_224_module_data_in[5] ,
    \sw_224_module_data_in[4] ,
    \sw_224_module_data_in[3] ,
    \sw_224_module_data_in[2] ,
    \sw_224_module_data_in[1] ,
    \sw_224_module_data_in[0] }),
    .module_data_out({\sw_224_module_data_out[7] ,
    \sw_224_module_data_out[6] ,
    \sw_224_module_data_out[5] ,
    \sw_224_module_data_out[4] ,
    \sw_224_module_data_out[3] ,
    \sw_224_module_data_out[2] ,
    \sw_224_module_data_out[1] ,
    \sw_224_module_data_out[0] }));
 scanchain scanchain_225 (.clk_in(sw_224_clk_out),
    .clk_out(sw_225_clk_out),
    .data_in(sw_224_data_out),
    .data_out(sw_225_data_out),
    .latch_enable_in(sw_224_latch_out),
    .latch_enable_out(sw_225_latch_out),
    .scan_select_in(sw_224_scan_out),
    .scan_select_out(sw_225_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_225_module_data_in[7] ,
    \sw_225_module_data_in[6] ,
    \sw_225_module_data_in[5] ,
    \sw_225_module_data_in[4] ,
    \sw_225_module_data_in[3] ,
    \sw_225_module_data_in[2] ,
    \sw_225_module_data_in[1] ,
    \sw_225_module_data_in[0] }),
    .module_data_out({\sw_225_module_data_out[7] ,
    \sw_225_module_data_out[6] ,
    \sw_225_module_data_out[5] ,
    \sw_225_module_data_out[4] ,
    \sw_225_module_data_out[3] ,
    \sw_225_module_data_out[2] ,
    \sw_225_module_data_out[1] ,
    \sw_225_module_data_out[0] }));
 scanchain scanchain_226 (.clk_in(sw_225_clk_out),
    .clk_out(sw_226_clk_out),
    .data_in(sw_225_data_out),
    .data_out(sw_226_data_out),
    .latch_enable_in(sw_225_latch_out),
    .latch_enable_out(sw_226_latch_out),
    .scan_select_in(sw_225_scan_out),
    .scan_select_out(sw_226_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_226_module_data_in[7] ,
    \sw_226_module_data_in[6] ,
    \sw_226_module_data_in[5] ,
    \sw_226_module_data_in[4] ,
    \sw_226_module_data_in[3] ,
    \sw_226_module_data_in[2] ,
    \sw_226_module_data_in[1] ,
    \sw_226_module_data_in[0] }),
    .module_data_out({\sw_226_module_data_out[7] ,
    \sw_226_module_data_out[6] ,
    \sw_226_module_data_out[5] ,
    \sw_226_module_data_out[4] ,
    \sw_226_module_data_out[3] ,
    \sw_226_module_data_out[2] ,
    \sw_226_module_data_out[1] ,
    \sw_226_module_data_out[0] }));
 scanchain scanchain_227 (.clk_in(sw_226_clk_out),
    .clk_out(sw_227_clk_out),
    .data_in(sw_226_data_out),
    .data_out(sw_227_data_out),
    .latch_enable_in(sw_226_latch_out),
    .latch_enable_out(sw_227_latch_out),
    .scan_select_in(sw_226_scan_out),
    .scan_select_out(sw_227_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_227_module_data_in[7] ,
    \sw_227_module_data_in[6] ,
    \sw_227_module_data_in[5] ,
    \sw_227_module_data_in[4] ,
    \sw_227_module_data_in[3] ,
    \sw_227_module_data_in[2] ,
    \sw_227_module_data_in[1] ,
    \sw_227_module_data_in[0] }),
    .module_data_out({\sw_227_module_data_out[7] ,
    \sw_227_module_data_out[6] ,
    \sw_227_module_data_out[5] ,
    \sw_227_module_data_out[4] ,
    \sw_227_module_data_out[3] ,
    \sw_227_module_data_out[2] ,
    \sw_227_module_data_out[1] ,
    \sw_227_module_data_out[0] }));
 scanchain scanchain_228 (.clk_in(sw_227_clk_out),
    .clk_out(sw_228_clk_out),
    .data_in(sw_227_data_out),
    .data_out(sw_228_data_out),
    .latch_enable_in(sw_227_latch_out),
    .latch_enable_out(sw_228_latch_out),
    .scan_select_in(sw_227_scan_out),
    .scan_select_out(sw_228_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_228_module_data_in[7] ,
    \sw_228_module_data_in[6] ,
    \sw_228_module_data_in[5] ,
    \sw_228_module_data_in[4] ,
    \sw_228_module_data_in[3] ,
    \sw_228_module_data_in[2] ,
    \sw_228_module_data_in[1] ,
    \sw_228_module_data_in[0] }),
    .module_data_out({\sw_228_module_data_out[7] ,
    \sw_228_module_data_out[6] ,
    \sw_228_module_data_out[5] ,
    \sw_228_module_data_out[4] ,
    \sw_228_module_data_out[3] ,
    \sw_228_module_data_out[2] ,
    \sw_228_module_data_out[1] ,
    \sw_228_module_data_out[0] }));
 scanchain scanchain_229 (.clk_in(sw_228_clk_out),
    .clk_out(sw_229_clk_out),
    .data_in(sw_228_data_out),
    .data_out(sw_229_data_out),
    .latch_enable_in(sw_228_latch_out),
    .latch_enable_out(sw_229_latch_out),
    .scan_select_in(sw_228_scan_out),
    .scan_select_out(sw_229_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_229_module_data_in[7] ,
    \sw_229_module_data_in[6] ,
    \sw_229_module_data_in[5] ,
    \sw_229_module_data_in[4] ,
    \sw_229_module_data_in[3] ,
    \sw_229_module_data_in[2] ,
    \sw_229_module_data_in[1] ,
    \sw_229_module_data_in[0] }),
    .module_data_out({\sw_229_module_data_out[7] ,
    \sw_229_module_data_out[6] ,
    \sw_229_module_data_out[5] ,
    \sw_229_module_data_out[4] ,
    \sw_229_module_data_out[3] ,
    \sw_229_module_data_out[2] ,
    \sw_229_module_data_out[1] ,
    \sw_229_module_data_out[0] }));
 scanchain scanchain_230 (.clk_in(sw_229_clk_out),
    .clk_out(sw_230_clk_out),
    .data_in(sw_229_data_out),
    .data_out(sw_230_data_out),
    .latch_enable_in(sw_229_latch_out),
    .latch_enable_out(sw_230_latch_out),
    .scan_select_in(sw_229_scan_out),
    .scan_select_out(sw_230_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_230_module_data_in[7] ,
    \sw_230_module_data_in[6] ,
    \sw_230_module_data_in[5] ,
    \sw_230_module_data_in[4] ,
    \sw_230_module_data_in[3] ,
    \sw_230_module_data_in[2] ,
    \sw_230_module_data_in[1] ,
    \sw_230_module_data_in[0] }),
    .module_data_out({\sw_230_module_data_out[7] ,
    \sw_230_module_data_out[6] ,
    \sw_230_module_data_out[5] ,
    \sw_230_module_data_out[4] ,
    \sw_230_module_data_out[3] ,
    \sw_230_module_data_out[2] ,
    \sw_230_module_data_out[1] ,
    \sw_230_module_data_out[0] }));
 scanchain scanchain_231 (.clk_in(sw_230_clk_out),
    .clk_out(sw_231_clk_out),
    .data_in(sw_230_data_out),
    .data_out(sw_231_data_out),
    .latch_enable_in(sw_230_latch_out),
    .latch_enable_out(sw_231_latch_out),
    .scan_select_in(sw_230_scan_out),
    .scan_select_out(sw_231_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_231_module_data_in[7] ,
    \sw_231_module_data_in[6] ,
    \sw_231_module_data_in[5] ,
    \sw_231_module_data_in[4] ,
    \sw_231_module_data_in[3] ,
    \sw_231_module_data_in[2] ,
    \sw_231_module_data_in[1] ,
    \sw_231_module_data_in[0] }),
    .module_data_out({\sw_231_module_data_out[7] ,
    \sw_231_module_data_out[6] ,
    \sw_231_module_data_out[5] ,
    \sw_231_module_data_out[4] ,
    \sw_231_module_data_out[3] ,
    \sw_231_module_data_out[2] ,
    \sw_231_module_data_out[1] ,
    \sw_231_module_data_out[0] }));
 scanchain scanchain_232 (.clk_in(sw_231_clk_out),
    .clk_out(sw_232_clk_out),
    .data_in(sw_231_data_out),
    .data_out(sw_232_data_out),
    .latch_enable_in(sw_231_latch_out),
    .latch_enable_out(sw_232_latch_out),
    .scan_select_in(sw_231_scan_out),
    .scan_select_out(sw_232_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_232_module_data_in[7] ,
    \sw_232_module_data_in[6] ,
    \sw_232_module_data_in[5] ,
    \sw_232_module_data_in[4] ,
    \sw_232_module_data_in[3] ,
    \sw_232_module_data_in[2] ,
    \sw_232_module_data_in[1] ,
    \sw_232_module_data_in[0] }),
    .module_data_out({\sw_232_module_data_out[7] ,
    \sw_232_module_data_out[6] ,
    \sw_232_module_data_out[5] ,
    \sw_232_module_data_out[4] ,
    \sw_232_module_data_out[3] ,
    \sw_232_module_data_out[2] ,
    \sw_232_module_data_out[1] ,
    \sw_232_module_data_out[0] }));
 scanchain scanchain_233 (.clk_in(sw_232_clk_out),
    .clk_out(sw_233_clk_out),
    .data_in(sw_232_data_out),
    .data_out(sw_233_data_out),
    .latch_enable_in(sw_232_latch_out),
    .latch_enable_out(sw_233_latch_out),
    .scan_select_in(sw_232_scan_out),
    .scan_select_out(sw_233_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_233_module_data_in[7] ,
    \sw_233_module_data_in[6] ,
    \sw_233_module_data_in[5] ,
    \sw_233_module_data_in[4] ,
    \sw_233_module_data_in[3] ,
    \sw_233_module_data_in[2] ,
    \sw_233_module_data_in[1] ,
    \sw_233_module_data_in[0] }),
    .module_data_out({\sw_233_module_data_out[7] ,
    \sw_233_module_data_out[6] ,
    \sw_233_module_data_out[5] ,
    \sw_233_module_data_out[4] ,
    \sw_233_module_data_out[3] ,
    \sw_233_module_data_out[2] ,
    \sw_233_module_data_out[1] ,
    \sw_233_module_data_out[0] }));
 scanchain scanchain_234 (.clk_in(sw_233_clk_out),
    .clk_out(sw_234_clk_out),
    .data_in(sw_233_data_out),
    .data_out(sw_234_data_out),
    .latch_enable_in(sw_233_latch_out),
    .latch_enable_out(sw_234_latch_out),
    .scan_select_in(sw_233_scan_out),
    .scan_select_out(sw_234_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_234_module_data_in[7] ,
    \sw_234_module_data_in[6] ,
    \sw_234_module_data_in[5] ,
    \sw_234_module_data_in[4] ,
    \sw_234_module_data_in[3] ,
    \sw_234_module_data_in[2] ,
    \sw_234_module_data_in[1] ,
    \sw_234_module_data_in[0] }),
    .module_data_out({\sw_234_module_data_out[7] ,
    \sw_234_module_data_out[6] ,
    \sw_234_module_data_out[5] ,
    \sw_234_module_data_out[4] ,
    \sw_234_module_data_out[3] ,
    \sw_234_module_data_out[2] ,
    \sw_234_module_data_out[1] ,
    \sw_234_module_data_out[0] }));
 scanchain scanchain_235 (.clk_in(sw_234_clk_out),
    .clk_out(sw_235_clk_out),
    .data_in(sw_234_data_out),
    .data_out(sw_235_data_out),
    .latch_enable_in(sw_234_latch_out),
    .latch_enable_out(sw_235_latch_out),
    .scan_select_in(sw_234_scan_out),
    .scan_select_out(sw_235_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_235_module_data_in[7] ,
    \sw_235_module_data_in[6] ,
    \sw_235_module_data_in[5] ,
    \sw_235_module_data_in[4] ,
    \sw_235_module_data_in[3] ,
    \sw_235_module_data_in[2] ,
    \sw_235_module_data_in[1] ,
    \sw_235_module_data_in[0] }),
    .module_data_out({\sw_235_module_data_out[7] ,
    \sw_235_module_data_out[6] ,
    \sw_235_module_data_out[5] ,
    \sw_235_module_data_out[4] ,
    \sw_235_module_data_out[3] ,
    \sw_235_module_data_out[2] ,
    \sw_235_module_data_out[1] ,
    \sw_235_module_data_out[0] }));
 scanchain scanchain_236 (.clk_in(sw_235_clk_out),
    .clk_out(sw_236_clk_out),
    .data_in(sw_235_data_out),
    .data_out(sw_236_data_out),
    .latch_enable_in(sw_235_latch_out),
    .latch_enable_out(sw_236_latch_out),
    .scan_select_in(sw_235_scan_out),
    .scan_select_out(sw_236_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_236_module_data_in[7] ,
    \sw_236_module_data_in[6] ,
    \sw_236_module_data_in[5] ,
    \sw_236_module_data_in[4] ,
    \sw_236_module_data_in[3] ,
    \sw_236_module_data_in[2] ,
    \sw_236_module_data_in[1] ,
    \sw_236_module_data_in[0] }),
    .module_data_out({\sw_236_module_data_out[7] ,
    \sw_236_module_data_out[6] ,
    \sw_236_module_data_out[5] ,
    \sw_236_module_data_out[4] ,
    \sw_236_module_data_out[3] ,
    \sw_236_module_data_out[2] ,
    \sw_236_module_data_out[1] ,
    \sw_236_module_data_out[0] }));
 scanchain scanchain_237 (.clk_in(sw_236_clk_out),
    .clk_out(sw_237_clk_out),
    .data_in(sw_236_data_out),
    .data_out(sw_237_data_out),
    .latch_enable_in(sw_236_latch_out),
    .latch_enable_out(sw_237_latch_out),
    .scan_select_in(sw_236_scan_out),
    .scan_select_out(sw_237_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_237_module_data_in[7] ,
    \sw_237_module_data_in[6] ,
    \sw_237_module_data_in[5] ,
    \sw_237_module_data_in[4] ,
    \sw_237_module_data_in[3] ,
    \sw_237_module_data_in[2] ,
    \sw_237_module_data_in[1] ,
    \sw_237_module_data_in[0] }),
    .module_data_out({\sw_237_module_data_out[7] ,
    \sw_237_module_data_out[6] ,
    \sw_237_module_data_out[5] ,
    \sw_237_module_data_out[4] ,
    \sw_237_module_data_out[3] ,
    \sw_237_module_data_out[2] ,
    \sw_237_module_data_out[1] ,
    \sw_237_module_data_out[0] }));
 scanchain scanchain_238 (.clk_in(sw_237_clk_out),
    .clk_out(sw_238_clk_out),
    .data_in(sw_237_data_out),
    .data_out(sw_238_data_out),
    .latch_enable_in(sw_237_latch_out),
    .latch_enable_out(sw_238_latch_out),
    .scan_select_in(sw_237_scan_out),
    .scan_select_out(sw_238_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_238_module_data_in[7] ,
    \sw_238_module_data_in[6] ,
    \sw_238_module_data_in[5] ,
    \sw_238_module_data_in[4] ,
    \sw_238_module_data_in[3] ,
    \sw_238_module_data_in[2] ,
    \sw_238_module_data_in[1] ,
    \sw_238_module_data_in[0] }),
    .module_data_out({\sw_238_module_data_out[7] ,
    \sw_238_module_data_out[6] ,
    \sw_238_module_data_out[5] ,
    \sw_238_module_data_out[4] ,
    \sw_238_module_data_out[3] ,
    \sw_238_module_data_out[2] ,
    \sw_238_module_data_out[1] ,
    \sw_238_module_data_out[0] }));
 scanchain scanchain_239 (.clk_in(sw_238_clk_out),
    .clk_out(sw_239_clk_out),
    .data_in(sw_238_data_out),
    .data_out(sw_239_data_out),
    .latch_enable_in(sw_238_latch_out),
    .latch_enable_out(sw_239_latch_out),
    .scan_select_in(sw_238_scan_out),
    .scan_select_out(sw_239_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_239_module_data_in[7] ,
    \sw_239_module_data_in[6] ,
    \sw_239_module_data_in[5] ,
    \sw_239_module_data_in[4] ,
    \sw_239_module_data_in[3] ,
    \sw_239_module_data_in[2] ,
    \sw_239_module_data_in[1] ,
    \sw_239_module_data_in[0] }),
    .module_data_out({\sw_239_module_data_out[7] ,
    \sw_239_module_data_out[6] ,
    \sw_239_module_data_out[5] ,
    \sw_239_module_data_out[4] ,
    \sw_239_module_data_out[3] ,
    \sw_239_module_data_out[2] ,
    \sw_239_module_data_out[1] ,
    \sw_239_module_data_out[0] }));
 scanchain scanchain_240 (.clk_in(sw_239_clk_out),
    .clk_out(sw_240_clk_out),
    .data_in(sw_239_data_out),
    .data_out(sw_240_data_out),
    .latch_enable_in(sw_239_latch_out),
    .latch_enable_out(sw_240_latch_out),
    .scan_select_in(sw_239_scan_out),
    .scan_select_out(sw_240_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_240_module_data_in[7] ,
    \sw_240_module_data_in[6] ,
    \sw_240_module_data_in[5] ,
    \sw_240_module_data_in[4] ,
    \sw_240_module_data_in[3] ,
    \sw_240_module_data_in[2] ,
    \sw_240_module_data_in[1] ,
    \sw_240_module_data_in[0] }),
    .module_data_out({\sw_240_module_data_out[7] ,
    \sw_240_module_data_out[6] ,
    \sw_240_module_data_out[5] ,
    \sw_240_module_data_out[4] ,
    \sw_240_module_data_out[3] ,
    \sw_240_module_data_out[2] ,
    \sw_240_module_data_out[1] ,
    \sw_240_module_data_out[0] }));
 scanchain scanchain_241 (.clk_in(sw_240_clk_out),
    .clk_out(sw_241_clk_out),
    .data_in(sw_240_data_out),
    .data_out(sw_241_data_out),
    .latch_enable_in(sw_240_latch_out),
    .latch_enable_out(sw_241_latch_out),
    .scan_select_in(sw_240_scan_out),
    .scan_select_out(sw_241_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_241_module_data_in[7] ,
    \sw_241_module_data_in[6] ,
    \sw_241_module_data_in[5] ,
    \sw_241_module_data_in[4] ,
    \sw_241_module_data_in[3] ,
    \sw_241_module_data_in[2] ,
    \sw_241_module_data_in[1] ,
    \sw_241_module_data_in[0] }),
    .module_data_out({\sw_241_module_data_out[7] ,
    \sw_241_module_data_out[6] ,
    \sw_241_module_data_out[5] ,
    \sw_241_module_data_out[4] ,
    \sw_241_module_data_out[3] ,
    \sw_241_module_data_out[2] ,
    \sw_241_module_data_out[1] ,
    \sw_241_module_data_out[0] }));
 scanchain scanchain_242 (.clk_in(sw_241_clk_out),
    .clk_out(sw_242_clk_out),
    .data_in(sw_241_data_out),
    .data_out(sw_242_data_out),
    .latch_enable_in(sw_241_latch_out),
    .latch_enable_out(sw_242_latch_out),
    .scan_select_in(sw_241_scan_out),
    .scan_select_out(sw_242_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_242_module_data_in[7] ,
    \sw_242_module_data_in[6] ,
    \sw_242_module_data_in[5] ,
    \sw_242_module_data_in[4] ,
    \sw_242_module_data_in[3] ,
    \sw_242_module_data_in[2] ,
    \sw_242_module_data_in[1] ,
    \sw_242_module_data_in[0] }),
    .module_data_out({\sw_242_module_data_out[7] ,
    \sw_242_module_data_out[6] ,
    \sw_242_module_data_out[5] ,
    \sw_242_module_data_out[4] ,
    \sw_242_module_data_out[3] ,
    \sw_242_module_data_out[2] ,
    \sw_242_module_data_out[1] ,
    \sw_242_module_data_out[0] }));
 scanchain scanchain_243 (.clk_in(sw_242_clk_out),
    .clk_out(sw_243_clk_out),
    .data_in(sw_242_data_out),
    .data_out(sw_243_data_out),
    .latch_enable_in(sw_242_latch_out),
    .latch_enable_out(sw_243_latch_out),
    .scan_select_in(sw_242_scan_out),
    .scan_select_out(sw_243_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_243_module_data_in[7] ,
    \sw_243_module_data_in[6] ,
    \sw_243_module_data_in[5] ,
    \sw_243_module_data_in[4] ,
    \sw_243_module_data_in[3] ,
    \sw_243_module_data_in[2] ,
    \sw_243_module_data_in[1] ,
    \sw_243_module_data_in[0] }),
    .module_data_out({\sw_243_module_data_out[7] ,
    \sw_243_module_data_out[6] ,
    \sw_243_module_data_out[5] ,
    \sw_243_module_data_out[4] ,
    \sw_243_module_data_out[3] ,
    \sw_243_module_data_out[2] ,
    \sw_243_module_data_out[1] ,
    \sw_243_module_data_out[0] }));
 scanchain scanchain_244 (.clk_in(sw_243_clk_out),
    .clk_out(sw_244_clk_out),
    .data_in(sw_243_data_out),
    .data_out(sw_244_data_out),
    .latch_enable_in(sw_243_latch_out),
    .latch_enable_out(sw_244_latch_out),
    .scan_select_in(sw_243_scan_out),
    .scan_select_out(sw_244_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_244_module_data_in[7] ,
    \sw_244_module_data_in[6] ,
    \sw_244_module_data_in[5] ,
    \sw_244_module_data_in[4] ,
    \sw_244_module_data_in[3] ,
    \sw_244_module_data_in[2] ,
    \sw_244_module_data_in[1] ,
    \sw_244_module_data_in[0] }),
    .module_data_out({\sw_244_module_data_out[7] ,
    \sw_244_module_data_out[6] ,
    \sw_244_module_data_out[5] ,
    \sw_244_module_data_out[4] ,
    \sw_244_module_data_out[3] ,
    \sw_244_module_data_out[2] ,
    \sw_244_module_data_out[1] ,
    \sw_244_module_data_out[0] }));
 scanchain scanchain_245 (.clk_in(sw_244_clk_out),
    .clk_out(sw_245_clk_out),
    .data_in(sw_244_data_out),
    .data_out(sw_245_data_out),
    .latch_enable_in(sw_244_latch_out),
    .latch_enable_out(sw_245_latch_out),
    .scan_select_in(sw_244_scan_out),
    .scan_select_out(sw_245_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_245_module_data_in[7] ,
    \sw_245_module_data_in[6] ,
    \sw_245_module_data_in[5] ,
    \sw_245_module_data_in[4] ,
    \sw_245_module_data_in[3] ,
    \sw_245_module_data_in[2] ,
    \sw_245_module_data_in[1] ,
    \sw_245_module_data_in[0] }),
    .module_data_out({\sw_245_module_data_out[7] ,
    \sw_245_module_data_out[6] ,
    \sw_245_module_data_out[5] ,
    \sw_245_module_data_out[4] ,
    \sw_245_module_data_out[3] ,
    \sw_245_module_data_out[2] ,
    \sw_245_module_data_out[1] ,
    \sw_245_module_data_out[0] }));
 scanchain scanchain_246 (.clk_in(sw_245_clk_out),
    .clk_out(sw_246_clk_out),
    .data_in(sw_245_data_out),
    .data_out(sw_246_data_out),
    .latch_enable_in(sw_245_latch_out),
    .latch_enable_out(sw_246_latch_out),
    .scan_select_in(sw_245_scan_out),
    .scan_select_out(sw_246_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_246_module_data_in[7] ,
    \sw_246_module_data_in[6] ,
    \sw_246_module_data_in[5] ,
    \sw_246_module_data_in[4] ,
    \sw_246_module_data_in[3] ,
    \sw_246_module_data_in[2] ,
    \sw_246_module_data_in[1] ,
    \sw_246_module_data_in[0] }),
    .module_data_out({\sw_246_module_data_out[7] ,
    \sw_246_module_data_out[6] ,
    \sw_246_module_data_out[5] ,
    \sw_246_module_data_out[4] ,
    \sw_246_module_data_out[3] ,
    \sw_246_module_data_out[2] ,
    \sw_246_module_data_out[1] ,
    \sw_246_module_data_out[0] }));
 scanchain scanchain_247 (.clk_in(sw_246_clk_out),
    .clk_out(sw_247_clk_out),
    .data_in(sw_246_data_out),
    .data_out(sw_247_data_out),
    .latch_enable_in(sw_246_latch_out),
    .latch_enable_out(sw_247_latch_out),
    .scan_select_in(sw_246_scan_out),
    .scan_select_out(sw_247_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_247_module_data_in[7] ,
    \sw_247_module_data_in[6] ,
    \sw_247_module_data_in[5] ,
    \sw_247_module_data_in[4] ,
    \sw_247_module_data_in[3] ,
    \sw_247_module_data_in[2] ,
    \sw_247_module_data_in[1] ,
    \sw_247_module_data_in[0] }),
    .module_data_out({\sw_247_module_data_out[7] ,
    \sw_247_module_data_out[6] ,
    \sw_247_module_data_out[5] ,
    \sw_247_module_data_out[4] ,
    \sw_247_module_data_out[3] ,
    \sw_247_module_data_out[2] ,
    \sw_247_module_data_out[1] ,
    \sw_247_module_data_out[0] }));
 scanchain scanchain_248 (.clk_in(sw_247_clk_out),
    .clk_out(sw_248_clk_out),
    .data_in(sw_247_data_out),
    .data_out(sw_248_data_out),
    .latch_enable_in(sw_247_latch_out),
    .latch_enable_out(sw_248_latch_out),
    .scan_select_in(sw_247_scan_out),
    .scan_select_out(sw_248_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_248_module_data_in[7] ,
    \sw_248_module_data_in[6] ,
    \sw_248_module_data_in[5] ,
    \sw_248_module_data_in[4] ,
    \sw_248_module_data_in[3] ,
    \sw_248_module_data_in[2] ,
    \sw_248_module_data_in[1] ,
    \sw_248_module_data_in[0] }),
    .module_data_out({\sw_248_module_data_out[7] ,
    \sw_248_module_data_out[6] ,
    \sw_248_module_data_out[5] ,
    \sw_248_module_data_out[4] ,
    \sw_248_module_data_out[3] ,
    \sw_248_module_data_out[2] ,
    \sw_248_module_data_out[1] ,
    \sw_248_module_data_out[0] }));
 scanchain scanchain_249 (.clk_in(sw_248_clk_out),
    .clk_out(sc_clk_in),
    .data_in(sw_248_data_out),
    .data_out(sc_data_in),
    .latch_enable_in(sw_248_latch_out),
    .latch_enable_out(sw_249_latch_out),
    .scan_select_in(sw_248_scan_out),
    .scan_select_out(sw_249_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_249_module_data_in[7] ,
    \sw_249_module_data_in[6] ,
    \sw_249_module_data_in[5] ,
    \sw_249_module_data_in[4] ,
    \sw_249_module_data_in[3] ,
    \sw_249_module_data_in[2] ,
    \sw_249_module_data_in[1] ,
    \sw_249_module_data_in[0] }),
    .module_data_out({\sw_249_module_data_out[7] ,
    \sw_249_module_data_out[6] ,
    \sw_249_module_data_out[5] ,
    \sw_249_module_data_out[4] ,
    \sw_249_module_data_out[3] ,
    \sw_249_module_data_out[2] ,
    \sw_249_module_data_out[1] ,
    \sw_249_module_data_out[0] }));
 secretFile secretFile_145 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_145_module_data_in[7] ,
    \sw_145_module_data_in[6] ,
    \sw_145_module_data_in[5] ,
    \sw_145_module_data_in[4] ,
    \sw_145_module_data_in[3] ,
    \sw_145_module_data_in[2] ,
    \sw_145_module_data_in[1] ,
    \sw_145_module_data_in[0] }),
    .io_out({\sw_145_module_data_out[7] ,
    \sw_145_module_data_out[6] ,
    \sw_145_module_data_out[5] ,
    \sw_145_module_data_out[4] ,
    \sw_145_module_data_out[3] ,
    \sw_145_module_data_out[2] ,
    \sw_145_module_data_out[1] ,
    \sw_145_module_data_out[0] }));
 seven_segment_seconds seven_segment_seconds_157 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_157_module_data_in[7] ,
    \sw_157_module_data_in[6] ,
    \sw_157_module_data_in[5] ,
    \sw_157_module_data_in[4] ,
    \sw_157_module_data_in[3] ,
    \sw_157_module_data_in[2] ,
    \sw_157_module_data_in[1] ,
    \sw_157_module_data_in[0] }),
    .io_out({\sw_157_module_data_out[7] ,
    \sw_157_module_data_out[6] ,
    \sw_157_module_data_out[5] ,
    \sw_157_module_data_out[4] ,
    \sw_157_module_data_out[3] ,
    \sw_157_module_data_out[2] ,
    \sw_157_module_data_out[1] ,
    \sw_157_module_data_out[0] }));
 shan1293_2bitalu shan1293_2bitalu_104 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_104_module_data_in[7] ,
    \sw_104_module_data_in[6] ,
    \sw_104_module_data_in[5] ,
    \sw_104_module_data_in[4] ,
    \sw_104_module_data_in[3] ,
    \sw_104_module_data_in[2] ,
    \sw_104_module_data_in[1] ,
    \sw_104_module_data_in[0] }),
    .io_out({\sw_104_module_data_out[7] ,
    \sw_104_module_data_out[6] ,
    \sw_104_module_data_out[5] ,
    \sw_104_module_data_out[4] ,
    \sw_104_module_data_out[3] ,
    \sw_104_module_data_out[2] ,
    \sw_104_module_data_out[1] ,
    \sw_104_module_data_out[0] }));
 skullart skullart_165 (.vssd1(vssd1),
    .vccd1(vccd1));
 sophialiCMU_math sophialiCMU_math_149 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_149_module_data_in[7] ,
    \sw_149_module_data_in[6] ,
    \sw_149_module_data_in[5] ,
    \sw_149_module_data_in[4] ,
    \sw_149_module_data_in[3] ,
    \sw_149_module_data_in[2] ,
    \sw_149_module_data_in[1] ,
    \sw_149_module_data_in[0] }),
    .io_out({\sw_149_module_data_out[7] ,
    \sw_149_module_data_out[6] ,
    \sw_149_module_data_out[5] ,
    \sw_149_module_data_out[4] ,
    \sw_149_module_data_out[3] ,
    \sw_149_module_data_out[2] ,
    \sw_149_module_data_out[1] ,
    \sw_149_module_data_out[0] }));
 stevenmburns_toplevel stevenmburns_toplevel_119 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_119_module_data_in[7] ,
    \sw_119_module_data_in[6] ,
    \sw_119_module_data_in[5] ,
    \sw_119_module_data_in[4] ,
    \sw_119_module_data_in[3] ,
    \sw_119_module_data_in[2] ,
    \sw_119_module_data_in[1] ,
    \sw_119_module_data_in[0] }),
    .io_out({\sw_119_module_data_out[7] ,
    \sw_119_module_data_out[6] ,
    \sw_119_module_data_out[5] ,
    \sw_119_module_data_out[4] ,
    \sw_119_module_data_out[3] ,
    \sw_119_module_data_out[2] ,
    \sw_119_module_data_out[1] ,
    \sw_119_module_data_out[0] }));
 swalense_top swalense_top_115 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_115_module_data_in[7] ,
    \sw_115_module_data_in[6] ,
    \sw_115_module_data_in[5] ,
    \sw_115_module_data_in[4] ,
    \sw_115_module_data_in[3] ,
    \sw_115_module_data_in[2] ,
    \sw_115_module_data_in[1] ,
    \sw_115_module_data_in[0] }),
    .io_out({\sw_115_module_data_out[7] ,
    \sw_115_module_data_out[6] ,
    \sw_115_module_data_out[5] ,
    \sw_115_module_data_out[4] ,
    \sw_115_module_data_out[3] ,
    \sw_115_module_data_out[2] ,
    \sw_115_module_data_out[1] ,
    \sw_115_module_data_out[0] }));
 thezoq2_yafpga thezoq2_yafpga_038 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_038_module_data_in[7] ,
    \sw_038_module_data_in[6] ,
    \sw_038_module_data_in[5] ,
    \sw_038_module_data_in[4] ,
    \sw_038_module_data_in[3] ,
    \sw_038_module_data_in[2] ,
    \sw_038_module_data_in[1] ,
    \sw_038_module_data_in[0] }),
    .io_out({\sw_038_module_data_out[7] ,
    \sw_038_module_data_out[6] ,
    \sw_038_module_data_out[5] ,
    \sw_038_module_data_out[4] ,
    \sw_038_module_data_out[3] ,
    \sw_038_module_data_out[2] ,
    \sw_038_module_data_out[1] ,
    \sw_038_module_data_out[0] }));
 tholin_avalonsemi_5401 tholin_avalonsemi_5401_014 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_014_module_data_in[7] ,
    \sw_014_module_data_in[6] ,
    \sw_014_module_data_in[5] ,
    \sw_014_module_data_in[4] ,
    \sw_014_module_data_in[3] ,
    \sw_014_module_data_in[2] ,
    \sw_014_module_data_in[1] ,
    \sw_014_module_data_in[0] }),
    .io_out({\sw_014_module_data_out[7] ,
    \sw_014_module_data_out[6] ,
    \sw_014_module_data_out[5] ,
    \sw_014_module_data_out[4] ,
    \sw_014_module_data_out[3] ,
    \sw_014_module_data_out[2] ,
    \sw_014_module_data_out[1] ,
    \sw_014_module_data_out[0] }));
 tholin_avalonsemi_tbb1143 tholin_avalonsemi_tbb1143_024 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_024_module_data_in[7] ,
    \sw_024_module_data_in[6] ,
    \sw_024_module_data_in[5] ,
    \sw_024_module_data_in[4] ,
    \sw_024_module_data_in[3] ,
    \sw_024_module_data_in[2] ,
    \sw_024_module_data_in[1] ,
    \sw_024_module_data_in[0] }),
    .io_out({\sw_024_module_data_out[7] ,
    \sw_024_module_data_out[6] ,
    \sw_024_module_data_out[5] ,
    \sw_024_module_data_out[4] ,
    \sw_024_module_data_out[3] ,
    \sw_024_module_data_out[2] ,
    \sw_024_module_data_out[1] ,
    \sw_024_module_data_out[0] }));
 thunderbird_taillight_ctrl thunderbird_taillight_ctrl_089 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_089_module_data_in[7] ,
    \sw_089_module_data_in[6] ,
    \sw_089_module_data_in[5] ,
    \sw_089_module_data_in[4] ,
    \sw_089_module_data_in[3] ,
    \sw_089_module_data_in[2] ,
    \sw_089_module_data_in[1] ,
    \sw_089_module_data_in[0] }),
    .io_out({\sw_089_module_data_out[7] ,
    \sw_089_module_data_out[6] ,
    \sw_089_module_data_out[5] ,
    \sw_089_module_data_out[4] ,
    \sw_089_module_data_out[3] ,
    \sw_089_module_data_out[2] ,
    \sw_089_module_data_out[1] ,
    \sw_089_module_data_out[0] }));
 tiny_fft tiny_fft_015 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_015_module_data_in[7] ,
    \sw_015_module_data_in[6] ,
    \sw_015_module_data_in[5] ,
    \sw_015_module_data_in[4] ,
    \sw_015_module_data_in[3] ,
    \sw_015_module_data_in[2] ,
    \sw_015_module_data_in[1] ,
    \sw_015_module_data_in[0] }),
    .io_out({\sw_015_module_data_out[7] ,
    \sw_015_module_data_out[6] ,
    \sw_015_module_data_out[5] ,
    \sw_015_module_data_out[4] ,
    \sw_015_module_data_out[3] ,
    \sw_015_module_data_out[2] ,
    \sw_015_module_data_out[1] ,
    \sw_015_module_data_out[0] }));
 tiny_kinda_pic tiny_kinda_pic_106 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_106_module_data_in[7] ,
    \sw_106_module_data_in[6] ,
    \sw_106_module_data_in[5] ,
    \sw_106_module_data_in[4] ,
    \sw_106_module_data_in[3] ,
    \sw_106_module_data_in[2] ,
    \sw_106_module_data_in[1] ,
    \sw_106_module_data_in[0] }),
    .io_out({\sw_106_module_data_out[7] ,
    \sw_106_module_data_out[6] ,
    \sw_106_module_data_out[5] ,
    \sw_106_module_data_out[4] ,
    \sw_106_module_data_out[3] ,
    \sw_106_module_data_out[2] ,
    \sw_106_module_data_out[1] ,
    \sw_106_module_data_out[0] }));
 tomkeddie_top_tto tomkeddie_top_tto_002 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_002_module_data_in[7] ,
    \sw_002_module_data_in[6] ,
    \sw_002_module_data_in[5] ,
    \sw_002_module_data_in[4] ,
    \sw_002_module_data_in[3] ,
    \sw_002_module_data_in[2] ,
    \sw_002_module_data_in[1] ,
    \sw_002_module_data_in[0] }),
    .io_out({\sw_002_module_data_out[7] ,
    \sw_002_module_data_out[6] ,
    \sw_002_module_data_out[5] ,
    \sw_002_module_data_out[4] ,
    \sw_002_module_data_out[3] ,
    \sw_002_module_data_out[2] ,
    \sw_002_module_data_out[1] ,
    \sw_002_module_data_out[0] }));
 tomkeddie_top_tto_a tomkeddie_top_tto_a_025 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_025_module_data_in[7] ,
    \sw_025_module_data_in[6] ,
    \sw_025_module_data_in[5] ,
    \sw_025_module_data_in[4] ,
    \sw_025_module_data_in[3] ,
    \sw_025_module_data_in[2] ,
    \sw_025_module_data_in[1] ,
    \sw_025_module_data_in[0] }),
    .io_out({\sw_025_module_data_out[7] ,
    \sw_025_module_data_out[6] ,
    \sw_025_module_data_out[5] ,
    \sw_025_module_data_out[4] ,
    \sw_025_module_data_out[3] ,
    \sw_025_module_data_out[2] ,
    \sw_025_module_data_out[1] ,
    \sw_025_module_data_out[0] }));
 tt2_tholin_diceroll tt2_tholin_diceroll_061 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_061_module_data_in[7] ,
    \sw_061_module_data_in[6] ,
    \sw_061_module_data_in[5] ,
    \sw_061_module_data_in[4] ,
    \sw_061_module_data_in[3] ,
    \sw_061_module_data_in[2] ,
    \sw_061_module_data_in[1] ,
    \sw_061_module_data_in[0] }),
    .io_out({\sw_061_module_data_out[7] ,
    \sw_061_module_data_out[6] ,
    \sw_061_module_data_out[5] ,
    \sw_061_module_data_out[4] ,
    \sw_061_module_data_out[3] ,
    \sw_061_module_data_out[2] ,
    \sw_061_module_data_out[1] ,
    \sw_061_module_data_out[0] }));
 tt2_tholin_multiplexed_counter tt2_tholin_multiplexed_counter_050 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_050_module_data_in[7] ,
    \sw_050_module_data_in[6] ,
    \sw_050_module_data_in[5] ,
    \sw_050_module_data_in[4] ,
    \sw_050_module_data_in[3] ,
    \sw_050_module_data_in[2] ,
    \sw_050_module_data_in[1] ,
    \sw_050_module_data_in[0] }),
    .io_out({\sw_050_module_data_out[7] ,
    \sw_050_module_data_out[6] ,
    \sw_050_module_data_out[5] ,
    \sw_050_module_data_out[4] ,
    \sw_050_module_data_out[3] ,
    \sw_050_module_data_out[2] ,
    \sw_050_module_data_out[1] ,
    \sw_050_module_data_out[0] }));
 tt2_tholin_multiplier tt2_tholin_multiplier_049 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_049_module_data_in[7] ,
    \sw_049_module_data_in[6] ,
    \sw_049_module_data_in[5] ,
    \sw_049_module_data_in[4] ,
    \sw_049_module_data_in[3] ,
    \sw_049_module_data_in[2] ,
    \sw_049_module_data_in[1] ,
    \sw_049_module_data_in[0] }),
    .io_out({\sw_049_module_data_out[7] ,
    \sw_049_module_data_out[6] ,
    \sw_049_module_data_out[5] ,
    \sw_049_module_data_out[4] ,
    \sw_049_module_data_out[3] ,
    \sw_049_module_data_out[2] ,
    \sw_049_module_data_out[1] ,
    \sw_049_module_data_out[0] }));
 tt2_tholin_namebadge tt2_tholin_namebadge_056 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_056_module_data_in[7] ,
    \sw_056_module_data_in[6] ,
    \sw_056_module_data_in[5] ,
    \sw_056_module_data_in[4] ,
    \sw_056_module_data_in[3] ,
    \sw_056_module_data_in[2] ,
    \sw_056_module_data_in[1] ,
    \sw_056_module_data_in[0] }),
    .io_out({\sw_056_module_data_out[7] ,
    \sw_056_module_data_out[6] ,
    \sw_056_module_data_out[5] ,
    \sw_056_module_data_out[4] ,
    \sw_056_module_data_out[3] ,
    \sw_056_module_data_out[2] ,
    \sw_056_module_data_out[1] ,
    \sw_056_module_data_out[0] }));
 tucanae47_gray_ctr6 tucanae47_gray_ctr6_155 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_155_module_data_in[7] ,
    \sw_155_module_data_in[6] ,
    \sw_155_module_data_in[5] ,
    \sw_155_module_data_in[4] ,
    \sw_155_module_data_in[3] ,
    \sw_155_module_data_in[2] ,
    \sw_155_module_data_in[1] ,
    \sw_155_module_data_in[0] }),
    .io_out({\sw_155_module_data_out[7] ,
    \sw_155_module_data_out[6] ,
    \sw_155_module_data_out[5] ,
    \sw_155_module_data_out[4] ,
    \sw_155_module_data_out[3] ,
    \sw_155_module_data_out[2] ,
    \sw_155_module_data_out[1] ,
    \sw_155_module_data_out[0] }));
 udxs_sqrt_top udxs_sqrt_top_067 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_067_module_data_in[7] ,
    \sw_067_module_data_in[6] ,
    \sw_067_module_data_in[5] ,
    \sw_067_module_data_in[4] ,
    \sw_067_module_data_in[3] ,
    \sw_067_module_data_in[2] ,
    \sw_067_module_data_in[1] ,
    \sw_067_module_data_in[0] }),
    .io_out({\sw_067_module_data_out[7] ,
    \sw_067_module_data_out[6] ,
    \sw_067_module_data_out[5] ,
    \sw_067_module_data_out[4] ,
    \sw_067_module_data_out[3] ,
    \sw_067_module_data_out[2] ,
    \sw_067_module_data_out[1] ,
    \sw_067_module_data_out[0] }));
 user_module_339688086163161683 user_module_339688086163161683_159 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_159_module_data_in[7] ,
    \sw_159_module_data_in[6] ,
    \sw_159_module_data_in[5] ,
    \sw_159_module_data_in[4] ,
    \sw_159_module_data_in[3] ,
    \sw_159_module_data_in[2] ,
    \sw_159_module_data_in[1] ,
    \sw_159_module_data_in[0] }),
    .io_out({\sw_159_module_data_out[7] ,
    \sw_159_module_data_out[6] ,
    \sw_159_module_data_out[5] ,
    \sw_159_module_data_out[4] ,
    \sw_159_module_data_out[3] ,
    \sw_159_module_data_out[2] ,
    \sw_159_module_data_out[1] ,
    \sw_159_module_data_out[0] }));
 user_module_340318610245288530 user_module_340318610245288530_081 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_081_module_data_in[7] ,
    \sw_081_module_data_in[6] ,
    \sw_081_module_data_in[5] ,
    \sw_081_module_data_in[4] ,
    \sw_081_module_data_in[3] ,
    \sw_081_module_data_in[2] ,
    \sw_081_module_data_in[1] ,
    \sw_081_module_data_in[0] }),
    .io_out({\sw_081_module_data_out[7] ,
    \sw_081_module_data_out[6] ,
    \sw_081_module_data_out[5] ,
    \sw_081_module_data_out[4] ,
    \sw_081_module_data_out[3] ,
    \sw_081_module_data_out[2] ,
    \sw_081_module_data_out[1] ,
    \sw_081_module_data_out[0] }));
 user_module_340805072482992722 user_module_340805072482992722_156 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_156_module_data_in[7] ,
    \sw_156_module_data_in[6] ,
    \sw_156_module_data_in[5] ,
    \sw_156_module_data_in[4] ,
    \sw_156_module_data_in[3] ,
    \sw_156_module_data_in[2] ,
    \sw_156_module_data_in[1] ,
    \sw_156_module_data_in[0] }),
    .io_out({\sw_156_module_data_out[7] ,
    \sw_156_module_data_out[6] ,
    \sw_156_module_data_out[5] ,
    \sw_156_module_data_out[4] ,
    \sw_156_module_data_out[3] ,
    \sw_156_module_data_out[2] ,
    \sw_156_module_data_out[1] ,
    \sw_156_module_data_out[0] }));
 user_module_341164910646919762 user_module_341164910646919762_069 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_069_module_data_in[7] ,
    \sw_069_module_data_in[6] ,
    \sw_069_module_data_in[5] ,
    \sw_069_module_data_in[4] ,
    \sw_069_module_data_in[3] ,
    \sw_069_module_data_in[2] ,
    \sw_069_module_data_in[1] ,
    \sw_069_module_data_in[0] }),
    .io_out({\sw_069_module_data_out[7] ,
    \sw_069_module_data_out[6] ,
    \sw_069_module_data_out[5] ,
    \sw_069_module_data_out[4] ,
    \sw_069_module_data_out[3] ,
    \sw_069_module_data_out[2] ,
    \sw_069_module_data_out[1] ,
    \sw_069_module_data_out[0] }));
 user_module_341178154799333971 user_module_341178154799333971_086 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_086_module_data_in[7] ,
    \sw_086_module_data_in[6] ,
    \sw_086_module_data_in[5] ,
    \sw_086_module_data_in[4] ,
    \sw_086_module_data_in[3] ,
    \sw_086_module_data_in[2] ,
    \sw_086_module_data_in[1] ,
    \sw_086_module_data_in[0] }),
    .io_out({\sw_086_module_data_out[7] ,
    \sw_086_module_data_out[6] ,
    \sw_086_module_data_out[5] ,
    \sw_086_module_data_out[4] ,
    \sw_086_module_data_out[3] ,
    \sw_086_module_data_out[2] ,
    \sw_086_module_data_out[1] ,
    \sw_086_module_data_out[0] }));
 user_module_341178481588044372 user_module_341178481588044372_123 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_123_module_data_in[7] ,
    \sw_123_module_data_in[6] ,
    \sw_123_module_data_in[5] ,
    \sw_123_module_data_in[4] ,
    \sw_123_module_data_in[3] ,
    \sw_123_module_data_in[2] ,
    \sw_123_module_data_in[1] ,
    \sw_123_module_data_in[0] }),
    .io_out({\sw_123_module_data_out[7] ,
    \sw_123_module_data_out[6] ,
    \sw_123_module_data_out[5] ,
    \sw_123_module_data_out[4] ,
    \sw_123_module_data_out[3] ,
    \sw_123_module_data_out[2] ,
    \sw_123_module_data_out[1] ,
    \sw_123_module_data_out[0] }));
 user_module_341277789473735250 user_module_341277789473735250_095 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_095_module_data_in[7] ,
    \sw_095_module_data_in[6] ,
    \sw_095_module_data_in[5] ,
    \sw_095_module_data_in[4] ,
    \sw_095_module_data_in[3] ,
    \sw_095_module_data_in[2] ,
    \sw_095_module_data_in[1] ,
    \sw_095_module_data_in[0] }),
    .io_out({\sw_095_module_data_out[7] ,
    \sw_095_module_data_out[6] ,
    \sw_095_module_data_out[5] ,
    \sw_095_module_data_out[4] ,
    \sw_095_module_data_out[3] ,
    \sw_095_module_data_out[2] ,
    \sw_095_module_data_out[1] ,
    \sw_095_module_data_out[0] }));
 user_module_341279123277087315 user_module_341279123277087315_103 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_103_module_data_in[7] ,
    \sw_103_module_data_in[6] ,
    \sw_103_module_data_in[5] ,
    \sw_103_module_data_in[4] ,
    \sw_103_module_data_in[3] ,
    \sw_103_module_data_in[2] ,
    \sw_103_module_data_in[1] ,
    \sw_103_module_data_in[0] }),
    .io_out({\sw_103_module_data_out[7] ,
    \sw_103_module_data_out[6] ,
    \sw_103_module_data_out[5] ,
    \sw_103_module_data_out[4] ,
    \sw_103_module_data_out[3] ,
    \sw_103_module_data_out[2] ,
    \sw_103_module_data_out[1] ,
    \sw_103_module_data_out[0] }));
 user_module_341353928049295956 user_module_341353928049295956_154 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_154_module_data_in[7] ,
    \sw_154_module_data_in[6] ,
    \sw_154_module_data_in[5] ,
    \sw_154_module_data_in[4] ,
    \sw_154_module_data_in[3] ,
    \sw_154_module_data_in[2] ,
    \sw_154_module_data_in[1] ,
    \sw_154_module_data_in[0] }),
    .io_out({\sw_154_module_data_out[7] ,
    \sw_154_module_data_out[6] ,
    \sw_154_module_data_out[5] ,
    \sw_154_module_data_out[4] ,
    \sw_154_module_data_out[3] ,
    \sw_154_module_data_out[2] ,
    \sw_154_module_data_out[1] ,
    \sw_154_module_data_out[0] }));
 user_module_341423712597181012 user_module_341423712597181012_094 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_094_module_data_in[7] ,
    \sw_094_module_data_in[6] ,
    \sw_094_module_data_in[5] ,
    \sw_094_module_data_in[4] ,
    \sw_094_module_data_in[3] ,
    \sw_094_module_data_in[2] ,
    \sw_094_module_data_in[1] ,
    \sw_094_module_data_in[0] }),
    .io_out({\sw_094_module_data_out[7] ,
    \sw_094_module_data_out[6] ,
    \sw_094_module_data_out[5] ,
    \sw_094_module_data_out[4] ,
    \sw_094_module_data_out[3] ,
    \sw_094_module_data_out[2] ,
    \sw_094_module_data_out[1] ,
    \sw_094_module_data_out[0] }));
 user_module_341432030163108435 user_module_341432030163108435_108 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_108_module_data_in[7] ,
    \sw_108_module_data_in[6] ,
    \sw_108_module_data_in[5] ,
    \sw_108_module_data_in[4] ,
    \sw_108_module_data_in[3] ,
    \sw_108_module_data_in[2] ,
    \sw_108_module_data_in[1] ,
    \sw_108_module_data_in[0] }),
    .io_out({\sw_108_module_data_out[7] ,
    \sw_108_module_data_out[6] ,
    \sw_108_module_data_out[5] ,
    \sw_108_module_data_out[4] ,
    \sw_108_module_data_out[3] ,
    \sw_108_module_data_out[2] ,
    \sw_108_module_data_out[1] ,
    \sw_108_module_data_out[0] }));
 user_module_341438392303616596 user_module_341438392303616596_141 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_141_module_data_in[7] ,
    \sw_141_module_data_in[6] ,
    \sw_141_module_data_in[5] ,
    \sw_141_module_data_in[4] ,
    \sw_141_module_data_in[3] ,
    \sw_141_module_data_in[2] ,
    \sw_141_module_data_in[1] ,
    \sw_141_module_data_in[0] }),
    .io_out({\sw_141_module_data_out[7] ,
    \sw_141_module_data_out[6] ,
    \sw_141_module_data_out[5] ,
    \sw_141_module_data_out[4] ,
    \sw_141_module_data_out[3] ,
    \sw_141_module_data_out[2] ,
    \sw_141_module_data_out[1] ,
    \sw_141_module_data_out[0] }));
 user_module_341490465660469844 user_module_341490465660469844_065 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_065_module_data_in[7] ,
    \sw_065_module_data_in[6] ,
    \sw_065_module_data_in[5] ,
    \sw_065_module_data_in[4] ,
    \sw_065_module_data_in[3] ,
    \sw_065_module_data_in[2] ,
    \sw_065_module_data_in[1] ,
    \sw_065_module_data_in[0] }),
    .io_out({\sw_065_module_data_out[7] ,
    \sw_065_module_data_out[6] ,
    \sw_065_module_data_out[5] ,
    \sw_065_module_data_out[4] ,
    \sw_065_module_data_out[3] ,
    \sw_065_module_data_out[2] ,
    \sw_065_module_data_out[1] ,
    \sw_065_module_data_out[0] }));
 user_module_341516949939814994 user_module_341516949939814994_048 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_048_module_data_in[7] ,
    \sw_048_module_data_in[6] ,
    \sw_048_module_data_in[5] ,
    \sw_048_module_data_in[4] ,
    \sw_048_module_data_in[3] ,
    \sw_048_module_data_in[2] ,
    \sw_048_module_data_in[1] ,
    \sw_048_module_data_in[0] }),
    .io_out({\sw_048_module_data_out[7] ,
    \sw_048_module_data_out[6] ,
    \sw_048_module_data_out[5] ,
    \sw_048_module_data_out[4] ,
    \sw_048_module_data_out[3] ,
    \sw_048_module_data_out[2] ,
    \sw_048_module_data_out[1] ,
    \sw_048_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_000 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_000_module_data_in[7] ,
    \sw_000_module_data_in[6] ,
    \sw_000_module_data_in[5] ,
    \sw_000_module_data_in[4] ,
    \sw_000_module_data_in[3] ,
    \sw_000_module_data_in[2] ,
    \sw_000_module_data_in[1] ,
    \sw_000_module_data_in[0] }),
    .io_out({\sw_000_module_data_out[7] ,
    \sw_000_module_data_out[6] ,
    \sw_000_module_data_out[5] ,
    \sw_000_module_data_out[4] ,
    \sw_000_module_data_out[3] ,
    \sw_000_module_data_out[2] ,
    \sw_000_module_data_out[1] ,
    \sw_000_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_166 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_166_module_data_in[7] ,
    \sw_166_module_data_in[6] ,
    \sw_166_module_data_in[5] ,
    \sw_166_module_data_in[4] ,
    \sw_166_module_data_in[3] ,
    \sw_166_module_data_in[2] ,
    \sw_166_module_data_in[1] ,
    \sw_166_module_data_in[0] }),
    .io_out({\sw_166_module_data_out[7] ,
    \sw_166_module_data_out[6] ,
    \sw_166_module_data_out[5] ,
    \sw_166_module_data_out[4] ,
    \sw_166_module_data_out[3] ,
    \sw_166_module_data_out[2] ,
    \sw_166_module_data_out[1] ,
    \sw_166_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_167 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_167_module_data_in[7] ,
    \sw_167_module_data_in[6] ,
    \sw_167_module_data_in[5] ,
    \sw_167_module_data_in[4] ,
    \sw_167_module_data_in[3] ,
    \sw_167_module_data_in[2] ,
    \sw_167_module_data_in[1] ,
    \sw_167_module_data_in[0] }),
    .io_out({\sw_167_module_data_out[7] ,
    \sw_167_module_data_out[6] ,
    \sw_167_module_data_out[5] ,
    \sw_167_module_data_out[4] ,
    \sw_167_module_data_out[3] ,
    \sw_167_module_data_out[2] ,
    \sw_167_module_data_out[1] ,
    \sw_167_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_168 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_168_module_data_in[7] ,
    \sw_168_module_data_in[6] ,
    \sw_168_module_data_in[5] ,
    \sw_168_module_data_in[4] ,
    \sw_168_module_data_in[3] ,
    \sw_168_module_data_in[2] ,
    \sw_168_module_data_in[1] ,
    \sw_168_module_data_in[0] }),
    .io_out({\sw_168_module_data_out[7] ,
    \sw_168_module_data_out[6] ,
    \sw_168_module_data_out[5] ,
    \sw_168_module_data_out[4] ,
    \sw_168_module_data_out[3] ,
    \sw_168_module_data_out[2] ,
    \sw_168_module_data_out[1] ,
    \sw_168_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_169 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_169_module_data_in[7] ,
    \sw_169_module_data_in[6] ,
    \sw_169_module_data_in[5] ,
    \sw_169_module_data_in[4] ,
    \sw_169_module_data_in[3] ,
    \sw_169_module_data_in[2] ,
    \sw_169_module_data_in[1] ,
    \sw_169_module_data_in[0] }),
    .io_out({\sw_169_module_data_out[7] ,
    \sw_169_module_data_out[6] ,
    \sw_169_module_data_out[5] ,
    \sw_169_module_data_out[4] ,
    \sw_169_module_data_out[3] ,
    \sw_169_module_data_out[2] ,
    \sw_169_module_data_out[1] ,
    \sw_169_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_170 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_170_module_data_in[7] ,
    \sw_170_module_data_in[6] ,
    \sw_170_module_data_in[5] ,
    \sw_170_module_data_in[4] ,
    \sw_170_module_data_in[3] ,
    \sw_170_module_data_in[2] ,
    \sw_170_module_data_in[1] ,
    \sw_170_module_data_in[0] }),
    .io_out({\sw_170_module_data_out[7] ,
    \sw_170_module_data_out[6] ,
    \sw_170_module_data_out[5] ,
    \sw_170_module_data_out[4] ,
    \sw_170_module_data_out[3] ,
    \sw_170_module_data_out[2] ,
    \sw_170_module_data_out[1] ,
    \sw_170_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_171 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_171_module_data_in[7] ,
    \sw_171_module_data_in[6] ,
    \sw_171_module_data_in[5] ,
    \sw_171_module_data_in[4] ,
    \sw_171_module_data_in[3] ,
    \sw_171_module_data_in[2] ,
    \sw_171_module_data_in[1] ,
    \sw_171_module_data_in[0] }),
    .io_out({\sw_171_module_data_out[7] ,
    \sw_171_module_data_out[6] ,
    \sw_171_module_data_out[5] ,
    \sw_171_module_data_out[4] ,
    \sw_171_module_data_out[3] ,
    \sw_171_module_data_out[2] ,
    \sw_171_module_data_out[1] ,
    \sw_171_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_172 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_172_module_data_in[7] ,
    \sw_172_module_data_in[6] ,
    \sw_172_module_data_in[5] ,
    \sw_172_module_data_in[4] ,
    \sw_172_module_data_in[3] ,
    \sw_172_module_data_in[2] ,
    \sw_172_module_data_in[1] ,
    \sw_172_module_data_in[0] }),
    .io_out({\sw_172_module_data_out[7] ,
    \sw_172_module_data_out[6] ,
    \sw_172_module_data_out[5] ,
    \sw_172_module_data_out[4] ,
    \sw_172_module_data_out[3] ,
    \sw_172_module_data_out[2] ,
    \sw_172_module_data_out[1] ,
    \sw_172_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_173 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_173_module_data_in[7] ,
    \sw_173_module_data_in[6] ,
    \sw_173_module_data_in[5] ,
    \sw_173_module_data_in[4] ,
    \sw_173_module_data_in[3] ,
    \sw_173_module_data_in[2] ,
    \sw_173_module_data_in[1] ,
    \sw_173_module_data_in[0] }),
    .io_out({\sw_173_module_data_out[7] ,
    \sw_173_module_data_out[6] ,
    \sw_173_module_data_out[5] ,
    \sw_173_module_data_out[4] ,
    \sw_173_module_data_out[3] ,
    \sw_173_module_data_out[2] ,
    \sw_173_module_data_out[1] ,
    \sw_173_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_174 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_174_module_data_in[7] ,
    \sw_174_module_data_in[6] ,
    \sw_174_module_data_in[5] ,
    \sw_174_module_data_in[4] ,
    \sw_174_module_data_in[3] ,
    \sw_174_module_data_in[2] ,
    \sw_174_module_data_in[1] ,
    \sw_174_module_data_in[0] }),
    .io_out({\sw_174_module_data_out[7] ,
    \sw_174_module_data_out[6] ,
    \sw_174_module_data_out[5] ,
    \sw_174_module_data_out[4] ,
    \sw_174_module_data_out[3] ,
    \sw_174_module_data_out[2] ,
    \sw_174_module_data_out[1] ,
    \sw_174_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_175 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_175_module_data_in[7] ,
    \sw_175_module_data_in[6] ,
    \sw_175_module_data_in[5] ,
    \sw_175_module_data_in[4] ,
    \sw_175_module_data_in[3] ,
    \sw_175_module_data_in[2] ,
    \sw_175_module_data_in[1] ,
    \sw_175_module_data_in[0] }),
    .io_out({\sw_175_module_data_out[7] ,
    \sw_175_module_data_out[6] ,
    \sw_175_module_data_out[5] ,
    \sw_175_module_data_out[4] ,
    \sw_175_module_data_out[3] ,
    \sw_175_module_data_out[2] ,
    \sw_175_module_data_out[1] ,
    \sw_175_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_176 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_176_module_data_in[7] ,
    \sw_176_module_data_in[6] ,
    \sw_176_module_data_in[5] ,
    \sw_176_module_data_in[4] ,
    \sw_176_module_data_in[3] ,
    \sw_176_module_data_in[2] ,
    \sw_176_module_data_in[1] ,
    \sw_176_module_data_in[0] }),
    .io_out({\sw_176_module_data_out[7] ,
    \sw_176_module_data_out[6] ,
    \sw_176_module_data_out[5] ,
    \sw_176_module_data_out[4] ,
    \sw_176_module_data_out[3] ,
    \sw_176_module_data_out[2] ,
    \sw_176_module_data_out[1] ,
    \sw_176_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_177 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_177_module_data_in[7] ,
    \sw_177_module_data_in[6] ,
    \sw_177_module_data_in[5] ,
    \sw_177_module_data_in[4] ,
    \sw_177_module_data_in[3] ,
    \sw_177_module_data_in[2] ,
    \sw_177_module_data_in[1] ,
    \sw_177_module_data_in[0] }),
    .io_out({\sw_177_module_data_out[7] ,
    \sw_177_module_data_out[6] ,
    \sw_177_module_data_out[5] ,
    \sw_177_module_data_out[4] ,
    \sw_177_module_data_out[3] ,
    \sw_177_module_data_out[2] ,
    \sw_177_module_data_out[1] ,
    \sw_177_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_178 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_178_module_data_in[7] ,
    \sw_178_module_data_in[6] ,
    \sw_178_module_data_in[5] ,
    \sw_178_module_data_in[4] ,
    \sw_178_module_data_in[3] ,
    \sw_178_module_data_in[2] ,
    \sw_178_module_data_in[1] ,
    \sw_178_module_data_in[0] }),
    .io_out({\sw_178_module_data_out[7] ,
    \sw_178_module_data_out[6] ,
    \sw_178_module_data_out[5] ,
    \sw_178_module_data_out[4] ,
    \sw_178_module_data_out[3] ,
    \sw_178_module_data_out[2] ,
    \sw_178_module_data_out[1] ,
    \sw_178_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_179 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_179_module_data_in[7] ,
    \sw_179_module_data_in[6] ,
    \sw_179_module_data_in[5] ,
    \sw_179_module_data_in[4] ,
    \sw_179_module_data_in[3] ,
    \sw_179_module_data_in[2] ,
    \sw_179_module_data_in[1] ,
    \sw_179_module_data_in[0] }),
    .io_out({\sw_179_module_data_out[7] ,
    \sw_179_module_data_out[6] ,
    \sw_179_module_data_out[5] ,
    \sw_179_module_data_out[4] ,
    \sw_179_module_data_out[3] ,
    \sw_179_module_data_out[2] ,
    \sw_179_module_data_out[1] ,
    \sw_179_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_180 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_180_module_data_in[7] ,
    \sw_180_module_data_in[6] ,
    \sw_180_module_data_in[5] ,
    \sw_180_module_data_in[4] ,
    \sw_180_module_data_in[3] ,
    \sw_180_module_data_in[2] ,
    \sw_180_module_data_in[1] ,
    \sw_180_module_data_in[0] }),
    .io_out({\sw_180_module_data_out[7] ,
    \sw_180_module_data_out[6] ,
    \sw_180_module_data_out[5] ,
    \sw_180_module_data_out[4] ,
    \sw_180_module_data_out[3] ,
    \sw_180_module_data_out[2] ,
    \sw_180_module_data_out[1] ,
    \sw_180_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_181 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_181_module_data_in[7] ,
    \sw_181_module_data_in[6] ,
    \sw_181_module_data_in[5] ,
    \sw_181_module_data_in[4] ,
    \sw_181_module_data_in[3] ,
    \sw_181_module_data_in[2] ,
    \sw_181_module_data_in[1] ,
    \sw_181_module_data_in[0] }),
    .io_out({\sw_181_module_data_out[7] ,
    \sw_181_module_data_out[6] ,
    \sw_181_module_data_out[5] ,
    \sw_181_module_data_out[4] ,
    \sw_181_module_data_out[3] ,
    \sw_181_module_data_out[2] ,
    \sw_181_module_data_out[1] ,
    \sw_181_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_182 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_182_module_data_in[7] ,
    \sw_182_module_data_in[6] ,
    \sw_182_module_data_in[5] ,
    \sw_182_module_data_in[4] ,
    \sw_182_module_data_in[3] ,
    \sw_182_module_data_in[2] ,
    \sw_182_module_data_in[1] ,
    \sw_182_module_data_in[0] }),
    .io_out({\sw_182_module_data_out[7] ,
    \sw_182_module_data_out[6] ,
    \sw_182_module_data_out[5] ,
    \sw_182_module_data_out[4] ,
    \sw_182_module_data_out[3] ,
    \sw_182_module_data_out[2] ,
    \sw_182_module_data_out[1] ,
    \sw_182_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_183 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_183_module_data_in[7] ,
    \sw_183_module_data_in[6] ,
    \sw_183_module_data_in[5] ,
    \sw_183_module_data_in[4] ,
    \sw_183_module_data_in[3] ,
    \sw_183_module_data_in[2] ,
    \sw_183_module_data_in[1] ,
    \sw_183_module_data_in[0] }),
    .io_out({\sw_183_module_data_out[7] ,
    \sw_183_module_data_out[6] ,
    \sw_183_module_data_out[5] ,
    \sw_183_module_data_out[4] ,
    \sw_183_module_data_out[3] ,
    \sw_183_module_data_out[2] ,
    \sw_183_module_data_out[1] ,
    \sw_183_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_184 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_184_module_data_in[7] ,
    \sw_184_module_data_in[6] ,
    \sw_184_module_data_in[5] ,
    \sw_184_module_data_in[4] ,
    \sw_184_module_data_in[3] ,
    \sw_184_module_data_in[2] ,
    \sw_184_module_data_in[1] ,
    \sw_184_module_data_in[0] }),
    .io_out({\sw_184_module_data_out[7] ,
    \sw_184_module_data_out[6] ,
    \sw_184_module_data_out[5] ,
    \sw_184_module_data_out[4] ,
    \sw_184_module_data_out[3] ,
    \sw_184_module_data_out[2] ,
    \sw_184_module_data_out[1] ,
    \sw_184_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_185 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_185_module_data_in[7] ,
    \sw_185_module_data_in[6] ,
    \sw_185_module_data_in[5] ,
    \sw_185_module_data_in[4] ,
    \sw_185_module_data_in[3] ,
    \sw_185_module_data_in[2] ,
    \sw_185_module_data_in[1] ,
    \sw_185_module_data_in[0] }),
    .io_out({\sw_185_module_data_out[7] ,
    \sw_185_module_data_out[6] ,
    \sw_185_module_data_out[5] ,
    \sw_185_module_data_out[4] ,
    \sw_185_module_data_out[3] ,
    \sw_185_module_data_out[2] ,
    \sw_185_module_data_out[1] ,
    \sw_185_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_186 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_186_module_data_in[7] ,
    \sw_186_module_data_in[6] ,
    \sw_186_module_data_in[5] ,
    \sw_186_module_data_in[4] ,
    \sw_186_module_data_in[3] ,
    \sw_186_module_data_in[2] ,
    \sw_186_module_data_in[1] ,
    \sw_186_module_data_in[0] }),
    .io_out({\sw_186_module_data_out[7] ,
    \sw_186_module_data_out[6] ,
    \sw_186_module_data_out[5] ,
    \sw_186_module_data_out[4] ,
    \sw_186_module_data_out[3] ,
    \sw_186_module_data_out[2] ,
    \sw_186_module_data_out[1] ,
    \sw_186_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_187 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_187_module_data_in[7] ,
    \sw_187_module_data_in[6] ,
    \sw_187_module_data_in[5] ,
    \sw_187_module_data_in[4] ,
    \sw_187_module_data_in[3] ,
    \sw_187_module_data_in[2] ,
    \sw_187_module_data_in[1] ,
    \sw_187_module_data_in[0] }),
    .io_out({\sw_187_module_data_out[7] ,
    \sw_187_module_data_out[6] ,
    \sw_187_module_data_out[5] ,
    \sw_187_module_data_out[4] ,
    \sw_187_module_data_out[3] ,
    \sw_187_module_data_out[2] ,
    \sw_187_module_data_out[1] ,
    \sw_187_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_188 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_188_module_data_in[7] ,
    \sw_188_module_data_in[6] ,
    \sw_188_module_data_in[5] ,
    \sw_188_module_data_in[4] ,
    \sw_188_module_data_in[3] ,
    \sw_188_module_data_in[2] ,
    \sw_188_module_data_in[1] ,
    \sw_188_module_data_in[0] }),
    .io_out({\sw_188_module_data_out[7] ,
    \sw_188_module_data_out[6] ,
    \sw_188_module_data_out[5] ,
    \sw_188_module_data_out[4] ,
    \sw_188_module_data_out[3] ,
    \sw_188_module_data_out[2] ,
    \sw_188_module_data_out[1] ,
    \sw_188_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_189 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_189_module_data_in[7] ,
    \sw_189_module_data_in[6] ,
    \sw_189_module_data_in[5] ,
    \sw_189_module_data_in[4] ,
    \sw_189_module_data_in[3] ,
    \sw_189_module_data_in[2] ,
    \sw_189_module_data_in[1] ,
    \sw_189_module_data_in[0] }),
    .io_out({\sw_189_module_data_out[7] ,
    \sw_189_module_data_out[6] ,
    \sw_189_module_data_out[5] ,
    \sw_189_module_data_out[4] ,
    \sw_189_module_data_out[3] ,
    \sw_189_module_data_out[2] ,
    \sw_189_module_data_out[1] ,
    \sw_189_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_190 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_190_module_data_in[7] ,
    \sw_190_module_data_in[6] ,
    \sw_190_module_data_in[5] ,
    \sw_190_module_data_in[4] ,
    \sw_190_module_data_in[3] ,
    \sw_190_module_data_in[2] ,
    \sw_190_module_data_in[1] ,
    \sw_190_module_data_in[0] }),
    .io_out({\sw_190_module_data_out[7] ,
    \sw_190_module_data_out[6] ,
    \sw_190_module_data_out[5] ,
    \sw_190_module_data_out[4] ,
    \sw_190_module_data_out[3] ,
    \sw_190_module_data_out[2] ,
    \sw_190_module_data_out[1] ,
    \sw_190_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_191 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_191_module_data_in[7] ,
    \sw_191_module_data_in[6] ,
    \sw_191_module_data_in[5] ,
    \sw_191_module_data_in[4] ,
    \sw_191_module_data_in[3] ,
    \sw_191_module_data_in[2] ,
    \sw_191_module_data_in[1] ,
    \sw_191_module_data_in[0] }),
    .io_out({\sw_191_module_data_out[7] ,
    \sw_191_module_data_out[6] ,
    \sw_191_module_data_out[5] ,
    \sw_191_module_data_out[4] ,
    \sw_191_module_data_out[3] ,
    \sw_191_module_data_out[2] ,
    \sw_191_module_data_out[1] ,
    \sw_191_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_192 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_192_module_data_in[7] ,
    \sw_192_module_data_in[6] ,
    \sw_192_module_data_in[5] ,
    \sw_192_module_data_in[4] ,
    \sw_192_module_data_in[3] ,
    \sw_192_module_data_in[2] ,
    \sw_192_module_data_in[1] ,
    \sw_192_module_data_in[0] }),
    .io_out({\sw_192_module_data_out[7] ,
    \sw_192_module_data_out[6] ,
    \sw_192_module_data_out[5] ,
    \sw_192_module_data_out[4] ,
    \sw_192_module_data_out[3] ,
    \sw_192_module_data_out[2] ,
    \sw_192_module_data_out[1] ,
    \sw_192_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_193 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_193_module_data_in[7] ,
    \sw_193_module_data_in[6] ,
    \sw_193_module_data_in[5] ,
    \sw_193_module_data_in[4] ,
    \sw_193_module_data_in[3] ,
    \sw_193_module_data_in[2] ,
    \sw_193_module_data_in[1] ,
    \sw_193_module_data_in[0] }),
    .io_out({\sw_193_module_data_out[7] ,
    \sw_193_module_data_out[6] ,
    \sw_193_module_data_out[5] ,
    \sw_193_module_data_out[4] ,
    \sw_193_module_data_out[3] ,
    \sw_193_module_data_out[2] ,
    \sw_193_module_data_out[1] ,
    \sw_193_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_194 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_194_module_data_in[7] ,
    \sw_194_module_data_in[6] ,
    \sw_194_module_data_in[5] ,
    \sw_194_module_data_in[4] ,
    \sw_194_module_data_in[3] ,
    \sw_194_module_data_in[2] ,
    \sw_194_module_data_in[1] ,
    \sw_194_module_data_in[0] }),
    .io_out({\sw_194_module_data_out[7] ,
    \sw_194_module_data_out[6] ,
    \sw_194_module_data_out[5] ,
    \sw_194_module_data_out[4] ,
    \sw_194_module_data_out[3] ,
    \sw_194_module_data_out[2] ,
    \sw_194_module_data_out[1] ,
    \sw_194_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_195 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_195_module_data_in[7] ,
    \sw_195_module_data_in[6] ,
    \sw_195_module_data_in[5] ,
    \sw_195_module_data_in[4] ,
    \sw_195_module_data_in[3] ,
    \sw_195_module_data_in[2] ,
    \sw_195_module_data_in[1] ,
    \sw_195_module_data_in[0] }),
    .io_out({\sw_195_module_data_out[7] ,
    \sw_195_module_data_out[6] ,
    \sw_195_module_data_out[5] ,
    \sw_195_module_data_out[4] ,
    \sw_195_module_data_out[3] ,
    \sw_195_module_data_out[2] ,
    \sw_195_module_data_out[1] ,
    \sw_195_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_196 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_196_module_data_in[7] ,
    \sw_196_module_data_in[6] ,
    \sw_196_module_data_in[5] ,
    \sw_196_module_data_in[4] ,
    \sw_196_module_data_in[3] ,
    \sw_196_module_data_in[2] ,
    \sw_196_module_data_in[1] ,
    \sw_196_module_data_in[0] }),
    .io_out({\sw_196_module_data_out[7] ,
    \sw_196_module_data_out[6] ,
    \sw_196_module_data_out[5] ,
    \sw_196_module_data_out[4] ,
    \sw_196_module_data_out[3] ,
    \sw_196_module_data_out[2] ,
    \sw_196_module_data_out[1] ,
    \sw_196_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_197 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_197_module_data_in[7] ,
    \sw_197_module_data_in[6] ,
    \sw_197_module_data_in[5] ,
    \sw_197_module_data_in[4] ,
    \sw_197_module_data_in[3] ,
    \sw_197_module_data_in[2] ,
    \sw_197_module_data_in[1] ,
    \sw_197_module_data_in[0] }),
    .io_out({\sw_197_module_data_out[7] ,
    \sw_197_module_data_out[6] ,
    \sw_197_module_data_out[5] ,
    \sw_197_module_data_out[4] ,
    \sw_197_module_data_out[3] ,
    \sw_197_module_data_out[2] ,
    \sw_197_module_data_out[1] ,
    \sw_197_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_198 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_198_module_data_in[7] ,
    \sw_198_module_data_in[6] ,
    \sw_198_module_data_in[5] ,
    \sw_198_module_data_in[4] ,
    \sw_198_module_data_in[3] ,
    \sw_198_module_data_in[2] ,
    \sw_198_module_data_in[1] ,
    \sw_198_module_data_in[0] }),
    .io_out({\sw_198_module_data_out[7] ,
    \sw_198_module_data_out[6] ,
    \sw_198_module_data_out[5] ,
    \sw_198_module_data_out[4] ,
    \sw_198_module_data_out[3] ,
    \sw_198_module_data_out[2] ,
    \sw_198_module_data_out[1] ,
    \sw_198_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_199 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_199_module_data_in[7] ,
    \sw_199_module_data_in[6] ,
    \sw_199_module_data_in[5] ,
    \sw_199_module_data_in[4] ,
    \sw_199_module_data_in[3] ,
    \sw_199_module_data_in[2] ,
    \sw_199_module_data_in[1] ,
    \sw_199_module_data_in[0] }),
    .io_out({\sw_199_module_data_out[7] ,
    \sw_199_module_data_out[6] ,
    \sw_199_module_data_out[5] ,
    \sw_199_module_data_out[4] ,
    \sw_199_module_data_out[3] ,
    \sw_199_module_data_out[2] ,
    \sw_199_module_data_out[1] ,
    \sw_199_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_200 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_200_module_data_in[7] ,
    \sw_200_module_data_in[6] ,
    \sw_200_module_data_in[5] ,
    \sw_200_module_data_in[4] ,
    \sw_200_module_data_in[3] ,
    \sw_200_module_data_in[2] ,
    \sw_200_module_data_in[1] ,
    \sw_200_module_data_in[0] }),
    .io_out({\sw_200_module_data_out[7] ,
    \sw_200_module_data_out[6] ,
    \sw_200_module_data_out[5] ,
    \sw_200_module_data_out[4] ,
    \sw_200_module_data_out[3] ,
    \sw_200_module_data_out[2] ,
    \sw_200_module_data_out[1] ,
    \sw_200_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_201 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_201_module_data_in[7] ,
    \sw_201_module_data_in[6] ,
    \sw_201_module_data_in[5] ,
    \sw_201_module_data_in[4] ,
    \sw_201_module_data_in[3] ,
    \sw_201_module_data_in[2] ,
    \sw_201_module_data_in[1] ,
    \sw_201_module_data_in[0] }),
    .io_out({\sw_201_module_data_out[7] ,
    \sw_201_module_data_out[6] ,
    \sw_201_module_data_out[5] ,
    \sw_201_module_data_out[4] ,
    \sw_201_module_data_out[3] ,
    \sw_201_module_data_out[2] ,
    \sw_201_module_data_out[1] ,
    \sw_201_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_202 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_202_module_data_in[7] ,
    \sw_202_module_data_in[6] ,
    \sw_202_module_data_in[5] ,
    \sw_202_module_data_in[4] ,
    \sw_202_module_data_in[3] ,
    \sw_202_module_data_in[2] ,
    \sw_202_module_data_in[1] ,
    \sw_202_module_data_in[0] }),
    .io_out({\sw_202_module_data_out[7] ,
    \sw_202_module_data_out[6] ,
    \sw_202_module_data_out[5] ,
    \sw_202_module_data_out[4] ,
    \sw_202_module_data_out[3] ,
    \sw_202_module_data_out[2] ,
    \sw_202_module_data_out[1] ,
    \sw_202_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_203 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_203_module_data_in[7] ,
    \sw_203_module_data_in[6] ,
    \sw_203_module_data_in[5] ,
    \sw_203_module_data_in[4] ,
    \sw_203_module_data_in[3] ,
    \sw_203_module_data_in[2] ,
    \sw_203_module_data_in[1] ,
    \sw_203_module_data_in[0] }),
    .io_out({\sw_203_module_data_out[7] ,
    \sw_203_module_data_out[6] ,
    \sw_203_module_data_out[5] ,
    \sw_203_module_data_out[4] ,
    \sw_203_module_data_out[3] ,
    \sw_203_module_data_out[2] ,
    \sw_203_module_data_out[1] ,
    \sw_203_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_204 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_204_module_data_in[7] ,
    \sw_204_module_data_in[6] ,
    \sw_204_module_data_in[5] ,
    \sw_204_module_data_in[4] ,
    \sw_204_module_data_in[3] ,
    \sw_204_module_data_in[2] ,
    \sw_204_module_data_in[1] ,
    \sw_204_module_data_in[0] }),
    .io_out({\sw_204_module_data_out[7] ,
    \sw_204_module_data_out[6] ,
    \sw_204_module_data_out[5] ,
    \sw_204_module_data_out[4] ,
    \sw_204_module_data_out[3] ,
    \sw_204_module_data_out[2] ,
    \sw_204_module_data_out[1] ,
    \sw_204_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_205 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_205_module_data_in[7] ,
    \sw_205_module_data_in[6] ,
    \sw_205_module_data_in[5] ,
    \sw_205_module_data_in[4] ,
    \sw_205_module_data_in[3] ,
    \sw_205_module_data_in[2] ,
    \sw_205_module_data_in[1] ,
    \sw_205_module_data_in[0] }),
    .io_out({\sw_205_module_data_out[7] ,
    \sw_205_module_data_out[6] ,
    \sw_205_module_data_out[5] ,
    \sw_205_module_data_out[4] ,
    \sw_205_module_data_out[3] ,
    \sw_205_module_data_out[2] ,
    \sw_205_module_data_out[1] ,
    \sw_205_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_206 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_206_module_data_in[7] ,
    \sw_206_module_data_in[6] ,
    \sw_206_module_data_in[5] ,
    \sw_206_module_data_in[4] ,
    \sw_206_module_data_in[3] ,
    \sw_206_module_data_in[2] ,
    \sw_206_module_data_in[1] ,
    \sw_206_module_data_in[0] }),
    .io_out({\sw_206_module_data_out[7] ,
    \sw_206_module_data_out[6] ,
    \sw_206_module_data_out[5] ,
    \sw_206_module_data_out[4] ,
    \sw_206_module_data_out[3] ,
    \sw_206_module_data_out[2] ,
    \sw_206_module_data_out[1] ,
    \sw_206_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_207 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_207_module_data_in[7] ,
    \sw_207_module_data_in[6] ,
    \sw_207_module_data_in[5] ,
    \sw_207_module_data_in[4] ,
    \sw_207_module_data_in[3] ,
    \sw_207_module_data_in[2] ,
    \sw_207_module_data_in[1] ,
    \sw_207_module_data_in[0] }),
    .io_out({\sw_207_module_data_out[7] ,
    \sw_207_module_data_out[6] ,
    \sw_207_module_data_out[5] ,
    \sw_207_module_data_out[4] ,
    \sw_207_module_data_out[3] ,
    \sw_207_module_data_out[2] ,
    \sw_207_module_data_out[1] ,
    \sw_207_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_208 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_208_module_data_in[7] ,
    \sw_208_module_data_in[6] ,
    \sw_208_module_data_in[5] ,
    \sw_208_module_data_in[4] ,
    \sw_208_module_data_in[3] ,
    \sw_208_module_data_in[2] ,
    \sw_208_module_data_in[1] ,
    \sw_208_module_data_in[0] }),
    .io_out({\sw_208_module_data_out[7] ,
    \sw_208_module_data_out[6] ,
    \sw_208_module_data_out[5] ,
    \sw_208_module_data_out[4] ,
    \sw_208_module_data_out[3] ,
    \sw_208_module_data_out[2] ,
    \sw_208_module_data_out[1] ,
    \sw_208_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_209 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_209_module_data_in[7] ,
    \sw_209_module_data_in[6] ,
    \sw_209_module_data_in[5] ,
    \sw_209_module_data_in[4] ,
    \sw_209_module_data_in[3] ,
    \sw_209_module_data_in[2] ,
    \sw_209_module_data_in[1] ,
    \sw_209_module_data_in[0] }),
    .io_out({\sw_209_module_data_out[7] ,
    \sw_209_module_data_out[6] ,
    \sw_209_module_data_out[5] ,
    \sw_209_module_data_out[4] ,
    \sw_209_module_data_out[3] ,
    \sw_209_module_data_out[2] ,
    \sw_209_module_data_out[1] ,
    \sw_209_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_210 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_210_module_data_in[7] ,
    \sw_210_module_data_in[6] ,
    \sw_210_module_data_in[5] ,
    \sw_210_module_data_in[4] ,
    \sw_210_module_data_in[3] ,
    \sw_210_module_data_in[2] ,
    \sw_210_module_data_in[1] ,
    \sw_210_module_data_in[0] }),
    .io_out({\sw_210_module_data_out[7] ,
    \sw_210_module_data_out[6] ,
    \sw_210_module_data_out[5] ,
    \sw_210_module_data_out[4] ,
    \sw_210_module_data_out[3] ,
    \sw_210_module_data_out[2] ,
    \sw_210_module_data_out[1] ,
    \sw_210_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_211 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_211_module_data_in[7] ,
    \sw_211_module_data_in[6] ,
    \sw_211_module_data_in[5] ,
    \sw_211_module_data_in[4] ,
    \sw_211_module_data_in[3] ,
    \sw_211_module_data_in[2] ,
    \sw_211_module_data_in[1] ,
    \sw_211_module_data_in[0] }),
    .io_out({\sw_211_module_data_out[7] ,
    \sw_211_module_data_out[6] ,
    \sw_211_module_data_out[5] ,
    \sw_211_module_data_out[4] ,
    \sw_211_module_data_out[3] ,
    \sw_211_module_data_out[2] ,
    \sw_211_module_data_out[1] ,
    \sw_211_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_212 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_212_module_data_in[7] ,
    \sw_212_module_data_in[6] ,
    \sw_212_module_data_in[5] ,
    \sw_212_module_data_in[4] ,
    \sw_212_module_data_in[3] ,
    \sw_212_module_data_in[2] ,
    \sw_212_module_data_in[1] ,
    \sw_212_module_data_in[0] }),
    .io_out({\sw_212_module_data_out[7] ,
    \sw_212_module_data_out[6] ,
    \sw_212_module_data_out[5] ,
    \sw_212_module_data_out[4] ,
    \sw_212_module_data_out[3] ,
    \sw_212_module_data_out[2] ,
    \sw_212_module_data_out[1] ,
    \sw_212_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_213 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_213_module_data_in[7] ,
    \sw_213_module_data_in[6] ,
    \sw_213_module_data_in[5] ,
    \sw_213_module_data_in[4] ,
    \sw_213_module_data_in[3] ,
    \sw_213_module_data_in[2] ,
    \sw_213_module_data_in[1] ,
    \sw_213_module_data_in[0] }),
    .io_out({\sw_213_module_data_out[7] ,
    \sw_213_module_data_out[6] ,
    \sw_213_module_data_out[5] ,
    \sw_213_module_data_out[4] ,
    \sw_213_module_data_out[3] ,
    \sw_213_module_data_out[2] ,
    \sw_213_module_data_out[1] ,
    \sw_213_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_214 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_214_module_data_in[7] ,
    \sw_214_module_data_in[6] ,
    \sw_214_module_data_in[5] ,
    \sw_214_module_data_in[4] ,
    \sw_214_module_data_in[3] ,
    \sw_214_module_data_in[2] ,
    \sw_214_module_data_in[1] ,
    \sw_214_module_data_in[0] }),
    .io_out({\sw_214_module_data_out[7] ,
    \sw_214_module_data_out[6] ,
    \sw_214_module_data_out[5] ,
    \sw_214_module_data_out[4] ,
    \sw_214_module_data_out[3] ,
    \sw_214_module_data_out[2] ,
    \sw_214_module_data_out[1] ,
    \sw_214_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_215 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_215_module_data_in[7] ,
    \sw_215_module_data_in[6] ,
    \sw_215_module_data_in[5] ,
    \sw_215_module_data_in[4] ,
    \sw_215_module_data_in[3] ,
    \sw_215_module_data_in[2] ,
    \sw_215_module_data_in[1] ,
    \sw_215_module_data_in[0] }),
    .io_out({\sw_215_module_data_out[7] ,
    \sw_215_module_data_out[6] ,
    \sw_215_module_data_out[5] ,
    \sw_215_module_data_out[4] ,
    \sw_215_module_data_out[3] ,
    \sw_215_module_data_out[2] ,
    \sw_215_module_data_out[1] ,
    \sw_215_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_216 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_216_module_data_in[7] ,
    \sw_216_module_data_in[6] ,
    \sw_216_module_data_in[5] ,
    \sw_216_module_data_in[4] ,
    \sw_216_module_data_in[3] ,
    \sw_216_module_data_in[2] ,
    \sw_216_module_data_in[1] ,
    \sw_216_module_data_in[0] }),
    .io_out({\sw_216_module_data_out[7] ,
    \sw_216_module_data_out[6] ,
    \sw_216_module_data_out[5] ,
    \sw_216_module_data_out[4] ,
    \sw_216_module_data_out[3] ,
    \sw_216_module_data_out[2] ,
    \sw_216_module_data_out[1] ,
    \sw_216_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_217 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_217_module_data_in[7] ,
    \sw_217_module_data_in[6] ,
    \sw_217_module_data_in[5] ,
    \sw_217_module_data_in[4] ,
    \sw_217_module_data_in[3] ,
    \sw_217_module_data_in[2] ,
    \sw_217_module_data_in[1] ,
    \sw_217_module_data_in[0] }),
    .io_out({\sw_217_module_data_out[7] ,
    \sw_217_module_data_out[6] ,
    \sw_217_module_data_out[5] ,
    \sw_217_module_data_out[4] ,
    \sw_217_module_data_out[3] ,
    \sw_217_module_data_out[2] ,
    \sw_217_module_data_out[1] ,
    \sw_217_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_218 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_218_module_data_in[7] ,
    \sw_218_module_data_in[6] ,
    \sw_218_module_data_in[5] ,
    \sw_218_module_data_in[4] ,
    \sw_218_module_data_in[3] ,
    \sw_218_module_data_in[2] ,
    \sw_218_module_data_in[1] ,
    \sw_218_module_data_in[0] }),
    .io_out({\sw_218_module_data_out[7] ,
    \sw_218_module_data_out[6] ,
    \sw_218_module_data_out[5] ,
    \sw_218_module_data_out[4] ,
    \sw_218_module_data_out[3] ,
    \sw_218_module_data_out[2] ,
    \sw_218_module_data_out[1] ,
    \sw_218_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_219 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_219_module_data_in[7] ,
    \sw_219_module_data_in[6] ,
    \sw_219_module_data_in[5] ,
    \sw_219_module_data_in[4] ,
    \sw_219_module_data_in[3] ,
    \sw_219_module_data_in[2] ,
    \sw_219_module_data_in[1] ,
    \sw_219_module_data_in[0] }),
    .io_out({\sw_219_module_data_out[7] ,
    \sw_219_module_data_out[6] ,
    \sw_219_module_data_out[5] ,
    \sw_219_module_data_out[4] ,
    \sw_219_module_data_out[3] ,
    \sw_219_module_data_out[2] ,
    \sw_219_module_data_out[1] ,
    \sw_219_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_220 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_220_module_data_in[7] ,
    \sw_220_module_data_in[6] ,
    \sw_220_module_data_in[5] ,
    \sw_220_module_data_in[4] ,
    \sw_220_module_data_in[3] ,
    \sw_220_module_data_in[2] ,
    \sw_220_module_data_in[1] ,
    \sw_220_module_data_in[0] }),
    .io_out({\sw_220_module_data_out[7] ,
    \sw_220_module_data_out[6] ,
    \sw_220_module_data_out[5] ,
    \sw_220_module_data_out[4] ,
    \sw_220_module_data_out[3] ,
    \sw_220_module_data_out[2] ,
    \sw_220_module_data_out[1] ,
    \sw_220_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_221 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_221_module_data_in[7] ,
    \sw_221_module_data_in[6] ,
    \sw_221_module_data_in[5] ,
    \sw_221_module_data_in[4] ,
    \sw_221_module_data_in[3] ,
    \sw_221_module_data_in[2] ,
    \sw_221_module_data_in[1] ,
    \sw_221_module_data_in[0] }),
    .io_out({\sw_221_module_data_out[7] ,
    \sw_221_module_data_out[6] ,
    \sw_221_module_data_out[5] ,
    \sw_221_module_data_out[4] ,
    \sw_221_module_data_out[3] ,
    \sw_221_module_data_out[2] ,
    \sw_221_module_data_out[1] ,
    \sw_221_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_222 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_222_module_data_in[7] ,
    \sw_222_module_data_in[6] ,
    \sw_222_module_data_in[5] ,
    \sw_222_module_data_in[4] ,
    \sw_222_module_data_in[3] ,
    \sw_222_module_data_in[2] ,
    \sw_222_module_data_in[1] ,
    \sw_222_module_data_in[0] }),
    .io_out({\sw_222_module_data_out[7] ,
    \sw_222_module_data_out[6] ,
    \sw_222_module_data_out[5] ,
    \sw_222_module_data_out[4] ,
    \sw_222_module_data_out[3] ,
    \sw_222_module_data_out[2] ,
    \sw_222_module_data_out[1] ,
    \sw_222_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_223 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_223_module_data_in[7] ,
    \sw_223_module_data_in[6] ,
    \sw_223_module_data_in[5] ,
    \sw_223_module_data_in[4] ,
    \sw_223_module_data_in[3] ,
    \sw_223_module_data_in[2] ,
    \sw_223_module_data_in[1] ,
    \sw_223_module_data_in[0] }),
    .io_out({\sw_223_module_data_out[7] ,
    \sw_223_module_data_out[6] ,
    \sw_223_module_data_out[5] ,
    \sw_223_module_data_out[4] ,
    \sw_223_module_data_out[3] ,
    \sw_223_module_data_out[2] ,
    \sw_223_module_data_out[1] ,
    \sw_223_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_224 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_224_module_data_in[7] ,
    \sw_224_module_data_in[6] ,
    \sw_224_module_data_in[5] ,
    \sw_224_module_data_in[4] ,
    \sw_224_module_data_in[3] ,
    \sw_224_module_data_in[2] ,
    \sw_224_module_data_in[1] ,
    \sw_224_module_data_in[0] }),
    .io_out({\sw_224_module_data_out[7] ,
    \sw_224_module_data_out[6] ,
    \sw_224_module_data_out[5] ,
    \sw_224_module_data_out[4] ,
    \sw_224_module_data_out[3] ,
    \sw_224_module_data_out[2] ,
    \sw_224_module_data_out[1] ,
    \sw_224_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_225 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_225_module_data_in[7] ,
    \sw_225_module_data_in[6] ,
    \sw_225_module_data_in[5] ,
    \sw_225_module_data_in[4] ,
    \sw_225_module_data_in[3] ,
    \sw_225_module_data_in[2] ,
    \sw_225_module_data_in[1] ,
    \sw_225_module_data_in[0] }),
    .io_out({\sw_225_module_data_out[7] ,
    \sw_225_module_data_out[6] ,
    \sw_225_module_data_out[5] ,
    \sw_225_module_data_out[4] ,
    \sw_225_module_data_out[3] ,
    \sw_225_module_data_out[2] ,
    \sw_225_module_data_out[1] ,
    \sw_225_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_226 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_226_module_data_in[7] ,
    \sw_226_module_data_in[6] ,
    \sw_226_module_data_in[5] ,
    \sw_226_module_data_in[4] ,
    \sw_226_module_data_in[3] ,
    \sw_226_module_data_in[2] ,
    \sw_226_module_data_in[1] ,
    \sw_226_module_data_in[0] }),
    .io_out({\sw_226_module_data_out[7] ,
    \sw_226_module_data_out[6] ,
    \sw_226_module_data_out[5] ,
    \sw_226_module_data_out[4] ,
    \sw_226_module_data_out[3] ,
    \sw_226_module_data_out[2] ,
    \sw_226_module_data_out[1] ,
    \sw_226_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_227 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_227_module_data_in[7] ,
    \sw_227_module_data_in[6] ,
    \sw_227_module_data_in[5] ,
    \sw_227_module_data_in[4] ,
    \sw_227_module_data_in[3] ,
    \sw_227_module_data_in[2] ,
    \sw_227_module_data_in[1] ,
    \sw_227_module_data_in[0] }),
    .io_out({\sw_227_module_data_out[7] ,
    \sw_227_module_data_out[6] ,
    \sw_227_module_data_out[5] ,
    \sw_227_module_data_out[4] ,
    \sw_227_module_data_out[3] ,
    \sw_227_module_data_out[2] ,
    \sw_227_module_data_out[1] ,
    \sw_227_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_228 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_228_module_data_in[7] ,
    \sw_228_module_data_in[6] ,
    \sw_228_module_data_in[5] ,
    \sw_228_module_data_in[4] ,
    \sw_228_module_data_in[3] ,
    \sw_228_module_data_in[2] ,
    \sw_228_module_data_in[1] ,
    \sw_228_module_data_in[0] }),
    .io_out({\sw_228_module_data_out[7] ,
    \sw_228_module_data_out[6] ,
    \sw_228_module_data_out[5] ,
    \sw_228_module_data_out[4] ,
    \sw_228_module_data_out[3] ,
    \sw_228_module_data_out[2] ,
    \sw_228_module_data_out[1] ,
    \sw_228_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_229 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_229_module_data_in[7] ,
    \sw_229_module_data_in[6] ,
    \sw_229_module_data_in[5] ,
    \sw_229_module_data_in[4] ,
    \sw_229_module_data_in[3] ,
    \sw_229_module_data_in[2] ,
    \sw_229_module_data_in[1] ,
    \sw_229_module_data_in[0] }),
    .io_out({\sw_229_module_data_out[7] ,
    \sw_229_module_data_out[6] ,
    \sw_229_module_data_out[5] ,
    \sw_229_module_data_out[4] ,
    \sw_229_module_data_out[3] ,
    \sw_229_module_data_out[2] ,
    \sw_229_module_data_out[1] ,
    \sw_229_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_230 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_230_module_data_in[7] ,
    \sw_230_module_data_in[6] ,
    \sw_230_module_data_in[5] ,
    \sw_230_module_data_in[4] ,
    \sw_230_module_data_in[3] ,
    \sw_230_module_data_in[2] ,
    \sw_230_module_data_in[1] ,
    \sw_230_module_data_in[0] }),
    .io_out({\sw_230_module_data_out[7] ,
    \sw_230_module_data_out[6] ,
    \sw_230_module_data_out[5] ,
    \sw_230_module_data_out[4] ,
    \sw_230_module_data_out[3] ,
    \sw_230_module_data_out[2] ,
    \sw_230_module_data_out[1] ,
    \sw_230_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_231 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_231_module_data_in[7] ,
    \sw_231_module_data_in[6] ,
    \sw_231_module_data_in[5] ,
    \sw_231_module_data_in[4] ,
    \sw_231_module_data_in[3] ,
    \sw_231_module_data_in[2] ,
    \sw_231_module_data_in[1] ,
    \sw_231_module_data_in[0] }),
    .io_out({\sw_231_module_data_out[7] ,
    \sw_231_module_data_out[6] ,
    \sw_231_module_data_out[5] ,
    \sw_231_module_data_out[4] ,
    \sw_231_module_data_out[3] ,
    \sw_231_module_data_out[2] ,
    \sw_231_module_data_out[1] ,
    \sw_231_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_232 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_232_module_data_in[7] ,
    \sw_232_module_data_in[6] ,
    \sw_232_module_data_in[5] ,
    \sw_232_module_data_in[4] ,
    \sw_232_module_data_in[3] ,
    \sw_232_module_data_in[2] ,
    \sw_232_module_data_in[1] ,
    \sw_232_module_data_in[0] }),
    .io_out({\sw_232_module_data_out[7] ,
    \sw_232_module_data_out[6] ,
    \sw_232_module_data_out[5] ,
    \sw_232_module_data_out[4] ,
    \sw_232_module_data_out[3] ,
    \sw_232_module_data_out[2] ,
    \sw_232_module_data_out[1] ,
    \sw_232_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_233 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_233_module_data_in[7] ,
    \sw_233_module_data_in[6] ,
    \sw_233_module_data_in[5] ,
    \sw_233_module_data_in[4] ,
    \sw_233_module_data_in[3] ,
    \sw_233_module_data_in[2] ,
    \sw_233_module_data_in[1] ,
    \sw_233_module_data_in[0] }),
    .io_out({\sw_233_module_data_out[7] ,
    \sw_233_module_data_out[6] ,
    \sw_233_module_data_out[5] ,
    \sw_233_module_data_out[4] ,
    \sw_233_module_data_out[3] ,
    \sw_233_module_data_out[2] ,
    \sw_233_module_data_out[1] ,
    \sw_233_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_234 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_234_module_data_in[7] ,
    \sw_234_module_data_in[6] ,
    \sw_234_module_data_in[5] ,
    \sw_234_module_data_in[4] ,
    \sw_234_module_data_in[3] ,
    \sw_234_module_data_in[2] ,
    \sw_234_module_data_in[1] ,
    \sw_234_module_data_in[0] }),
    .io_out({\sw_234_module_data_out[7] ,
    \sw_234_module_data_out[6] ,
    \sw_234_module_data_out[5] ,
    \sw_234_module_data_out[4] ,
    \sw_234_module_data_out[3] ,
    \sw_234_module_data_out[2] ,
    \sw_234_module_data_out[1] ,
    \sw_234_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_235 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_235_module_data_in[7] ,
    \sw_235_module_data_in[6] ,
    \sw_235_module_data_in[5] ,
    \sw_235_module_data_in[4] ,
    \sw_235_module_data_in[3] ,
    \sw_235_module_data_in[2] ,
    \sw_235_module_data_in[1] ,
    \sw_235_module_data_in[0] }),
    .io_out({\sw_235_module_data_out[7] ,
    \sw_235_module_data_out[6] ,
    \sw_235_module_data_out[5] ,
    \sw_235_module_data_out[4] ,
    \sw_235_module_data_out[3] ,
    \sw_235_module_data_out[2] ,
    \sw_235_module_data_out[1] ,
    \sw_235_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_236 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_236_module_data_in[7] ,
    \sw_236_module_data_in[6] ,
    \sw_236_module_data_in[5] ,
    \sw_236_module_data_in[4] ,
    \sw_236_module_data_in[3] ,
    \sw_236_module_data_in[2] ,
    \sw_236_module_data_in[1] ,
    \sw_236_module_data_in[0] }),
    .io_out({\sw_236_module_data_out[7] ,
    \sw_236_module_data_out[6] ,
    \sw_236_module_data_out[5] ,
    \sw_236_module_data_out[4] ,
    \sw_236_module_data_out[3] ,
    \sw_236_module_data_out[2] ,
    \sw_236_module_data_out[1] ,
    \sw_236_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_237 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_237_module_data_in[7] ,
    \sw_237_module_data_in[6] ,
    \sw_237_module_data_in[5] ,
    \sw_237_module_data_in[4] ,
    \sw_237_module_data_in[3] ,
    \sw_237_module_data_in[2] ,
    \sw_237_module_data_in[1] ,
    \sw_237_module_data_in[0] }),
    .io_out({\sw_237_module_data_out[7] ,
    \sw_237_module_data_out[6] ,
    \sw_237_module_data_out[5] ,
    \sw_237_module_data_out[4] ,
    \sw_237_module_data_out[3] ,
    \sw_237_module_data_out[2] ,
    \sw_237_module_data_out[1] ,
    \sw_237_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_238 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_238_module_data_in[7] ,
    \sw_238_module_data_in[6] ,
    \sw_238_module_data_in[5] ,
    \sw_238_module_data_in[4] ,
    \sw_238_module_data_in[3] ,
    \sw_238_module_data_in[2] ,
    \sw_238_module_data_in[1] ,
    \sw_238_module_data_in[0] }),
    .io_out({\sw_238_module_data_out[7] ,
    \sw_238_module_data_out[6] ,
    \sw_238_module_data_out[5] ,
    \sw_238_module_data_out[4] ,
    \sw_238_module_data_out[3] ,
    \sw_238_module_data_out[2] ,
    \sw_238_module_data_out[1] ,
    \sw_238_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_239 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_239_module_data_in[7] ,
    \sw_239_module_data_in[6] ,
    \sw_239_module_data_in[5] ,
    \sw_239_module_data_in[4] ,
    \sw_239_module_data_in[3] ,
    \sw_239_module_data_in[2] ,
    \sw_239_module_data_in[1] ,
    \sw_239_module_data_in[0] }),
    .io_out({\sw_239_module_data_out[7] ,
    \sw_239_module_data_out[6] ,
    \sw_239_module_data_out[5] ,
    \sw_239_module_data_out[4] ,
    \sw_239_module_data_out[3] ,
    \sw_239_module_data_out[2] ,
    \sw_239_module_data_out[1] ,
    \sw_239_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_240 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_240_module_data_in[7] ,
    \sw_240_module_data_in[6] ,
    \sw_240_module_data_in[5] ,
    \sw_240_module_data_in[4] ,
    \sw_240_module_data_in[3] ,
    \sw_240_module_data_in[2] ,
    \sw_240_module_data_in[1] ,
    \sw_240_module_data_in[0] }),
    .io_out({\sw_240_module_data_out[7] ,
    \sw_240_module_data_out[6] ,
    \sw_240_module_data_out[5] ,
    \sw_240_module_data_out[4] ,
    \sw_240_module_data_out[3] ,
    \sw_240_module_data_out[2] ,
    \sw_240_module_data_out[1] ,
    \sw_240_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_241 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_241_module_data_in[7] ,
    \sw_241_module_data_in[6] ,
    \sw_241_module_data_in[5] ,
    \sw_241_module_data_in[4] ,
    \sw_241_module_data_in[3] ,
    \sw_241_module_data_in[2] ,
    \sw_241_module_data_in[1] ,
    \sw_241_module_data_in[0] }),
    .io_out({\sw_241_module_data_out[7] ,
    \sw_241_module_data_out[6] ,
    \sw_241_module_data_out[5] ,
    \sw_241_module_data_out[4] ,
    \sw_241_module_data_out[3] ,
    \sw_241_module_data_out[2] ,
    \sw_241_module_data_out[1] ,
    \sw_241_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_242 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_242_module_data_in[7] ,
    \sw_242_module_data_in[6] ,
    \sw_242_module_data_in[5] ,
    \sw_242_module_data_in[4] ,
    \sw_242_module_data_in[3] ,
    \sw_242_module_data_in[2] ,
    \sw_242_module_data_in[1] ,
    \sw_242_module_data_in[0] }),
    .io_out({\sw_242_module_data_out[7] ,
    \sw_242_module_data_out[6] ,
    \sw_242_module_data_out[5] ,
    \sw_242_module_data_out[4] ,
    \sw_242_module_data_out[3] ,
    \sw_242_module_data_out[2] ,
    \sw_242_module_data_out[1] ,
    \sw_242_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_243 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_243_module_data_in[7] ,
    \sw_243_module_data_in[6] ,
    \sw_243_module_data_in[5] ,
    \sw_243_module_data_in[4] ,
    \sw_243_module_data_in[3] ,
    \sw_243_module_data_in[2] ,
    \sw_243_module_data_in[1] ,
    \sw_243_module_data_in[0] }),
    .io_out({\sw_243_module_data_out[7] ,
    \sw_243_module_data_out[6] ,
    \sw_243_module_data_out[5] ,
    \sw_243_module_data_out[4] ,
    \sw_243_module_data_out[3] ,
    \sw_243_module_data_out[2] ,
    \sw_243_module_data_out[1] ,
    \sw_243_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_244 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_244_module_data_in[7] ,
    \sw_244_module_data_in[6] ,
    \sw_244_module_data_in[5] ,
    \sw_244_module_data_in[4] ,
    \sw_244_module_data_in[3] ,
    \sw_244_module_data_in[2] ,
    \sw_244_module_data_in[1] ,
    \sw_244_module_data_in[0] }),
    .io_out({\sw_244_module_data_out[7] ,
    \sw_244_module_data_out[6] ,
    \sw_244_module_data_out[5] ,
    \sw_244_module_data_out[4] ,
    \sw_244_module_data_out[3] ,
    \sw_244_module_data_out[2] ,
    \sw_244_module_data_out[1] ,
    \sw_244_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_245 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_245_module_data_in[7] ,
    \sw_245_module_data_in[6] ,
    \sw_245_module_data_in[5] ,
    \sw_245_module_data_in[4] ,
    \sw_245_module_data_in[3] ,
    \sw_245_module_data_in[2] ,
    \sw_245_module_data_in[1] ,
    \sw_245_module_data_in[0] }),
    .io_out({\sw_245_module_data_out[7] ,
    \sw_245_module_data_out[6] ,
    \sw_245_module_data_out[5] ,
    \sw_245_module_data_out[4] ,
    \sw_245_module_data_out[3] ,
    \sw_245_module_data_out[2] ,
    \sw_245_module_data_out[1] ,
    \sw_245_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_246 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_246_module_data_in[7] ,
    \sw_246_module_data_in[6] ,
    \sw_246_module_data_in[5] ,
    \sw_246_module_data_in[4] ,
    \sw_246_module_data_in[3] ,
    \sw_246_module_data_in[2] ,
    \sw_246_module_data_in[1] ,
    \sw_246_module_data_in[0] }),
    .io_out({\sw_246_module_data_out[7] ,
    \sw_246_module_data_out[6] ,
    \sw_246_module_data_out[5] ,
    \sw_246_module_data_out[4] ,
    \sw_246_module_data_out[3] ,
    \sw_246_module_data_out[2] ,
    \sw_246_module_data_out[1] ,
    \sw_246_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_247 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_247_module_data_in[7] ,
    \sw_247_module_data_in[6] ,
    \sw_247_module_data_in[5] ,
    \sw_247_module_data_in[4] ,
    \sw_247_module_data_in[3] ,
    \sw_247_module_data_in[2] ,
    \sw_247_module_data_in[1] ,
    \sw_247_module_data_in[0] }),
    .io_out({\sw_247_module_data_out[7] ,
    \sw_247_module_data_out[6] ,
    \sw_247_module_data_out[5] ,
    \sw_247_module_data_out[4] ,
    \sw_247_module_data_out[3] ,
    \sw_247_module_data_out[2] ,
    \sw_247_module_data_out[1] ,
    \sw_247_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_248 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_248_module_data_in[7] ,
    \sw_248_module_data_in[6] ,
    \sw_248_module_data_in[5] ,
    \sw_248_module_data_in[4] ,
    \sw_248_module_data_in[3] ,
    \sw_248_module_data_in[2] ,
    \sw_248_module_data_in[1] ,
    \sw_248_module_data_in[0] }),
    .io_out({\sw_248_module_data_out[7] ,
    \sw_248_module_data_out[6] ,
    \sw_248_module_data_out[5] ,
    \sw_248_module_data_out[4] ,
    \sw_248_module_data_out[3] ,
    \sw_248_module_data_out[2] ,
    \sw_248_module_data_out[1] ,
    \sw_248_module_data_out[0] }));
 user_module_341535056611770964 user_module_341535056611770964_249 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_249_module_data_in[7] ,
    \sw_249_module_data_in[6] ,
    \sw_249_module_data_in[5] ,
    \sw_249_module_data_in[4] ,
    \sw_249_module_data_in[3] ,
    \sw_249_module_data_in[2] ,
    \sw_249_module_data_in[1] ,
    \sw_249_module_data_in[0] }),
    .io_out({\sw_249_module_data_out[7] ,
    \sw_249_module_data_out[6] ,
    \sw_249_module_data_out[5] ,
    \sw_249_module_data_out[4] ,
    \sw_249_module_data_out[3] ,
    \sw_249_module_data_out[2] ,
    \sw_249_module_data_out[1] ,
    \sw_249_module_data_out[0] }));
 user_module_341541108650607187 user_module_341541108650607187_047 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_047_module_data_in[7] ,
    \sw_047_module_data_in[6] ,
    \sw_047_module_data_in[5] ,
    \sw_047_module_data_in[4] ,
    \sw_047_module_data_in[3] ,
    \sw_047_module_data_in[2] ,
    \sw_047_module_data_in[1] ,
    \sw_047_module_data_in[0] }),
    .io_out({\sw_047_module_data_out[7] ,
    \sw_047_module_data_out[6] ,
    \sw_047_module_data_out[5] ,
    \sw_047_module_data_out[4] ,
    \sw_047_module_data_out[3] ,
    \sw_047_module_data_out[2] ,
    \sw_047_module_data_out[1] ,
    \sw_047_module_data_out[0] }));
 user_module_341546888233747026 user_module_341546888233747026_120 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_120_module_data_in[7] ,
    \sw_120_module_data_in[6] ,
    \sw_120_module_data_in[5] ,
    \sw_120_module_data_in[4] ,
    \sw_120_module_data_in[3] ,
    \sw_120_module_data_in[2] ,
    \sw_120_module_data_in[1] ,
    \sw_120_module_data_in[0] }),
    .io_out({\sw_120_module_data_out[7] ,
    \sw_120_module_data_out[6] ,
    \sw_120_module_data_out[5] ,
    \sw_120_module_data_out[4] ,
    \sw_120_module_data_out[3] ,
    \sw_120_module_data_out[2] ,
    \sw_120_module_data_out[1] ,
    \sw_120_module_data_out[0] }));
 user_module_341557831870186068 user_module_341557831870186068_140 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_140_module_data_in[7] ,
    \sw_140_module_data_in[6] ,
    \sw_140_module_data_in[5] ,
    \sw_140_module_data_in[4] ,
    \sw_140_module_data_in[3] ,
    \sw_140_module_data_in[2] ,
    \sw_140_module_data_in[1] ,
    \sw_140_module_data_in[0] }),
    .io_out({\sw_140_module_data_out[7] ,
    \sw_140_module_data_out[6] ,
    \sw_140_module_data_out[5] ,
    \sw_140_module_data_out[4] ,
    \sw_140_module_data_out[3] ,
    \sw_140_module_data_out[2] ,
    \sw_140_module_data_out[1] ,
    \sw_140_module_data_out[0] }));
 user_module_341571228858843732 user_module_341571228858843732_083 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_083_module_data_in[7] ,
    \sw_083_module_data_in[6] ,
    \sw_083_module_data_in[5] ,
    \sw_083_module_data_in[4] ,
    \sw_083_module_data_in[3] ,
    \sw_083_module_data_in[2] ,
    \sw_083_module_data_in[1] ,
    \sw_083_module_data_in[0] }),
    .io_out({\sw_083_module_data_out[7] ,
    \sw_083_module_data_out[6] ,
    \sw_083_module_data_out[5] ,
    \sw_083_module_data_out[4] ,
    \sw_083_module_data_out[3] ,
    \sw_083_module_data_out[2] ,
    \sw_083_module_data_out[1] ,
    \sw_083_module_data_out[0] }));
 user_module_341589685194195540 user_module_341589685194195540_091 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_091_module_data_in[7] ,
    \sw_091_module_data_in[6] ,
    \sw_091_module_data_in[5] ,
    \sw_091_module_data_in[4] ,
    \sw_091_module_data_in[3] ,
    \sw_091_module_data_in[2] ,
    \sw_091_module_data_in[1] ,
    \sw_091_module_data_in[0] }),
    .io_out({\sw_091_module_data_out[7] ,
    \sw_091_module_data_out[6] ,
    \sw_091_module_data_out[5] ,
    \sw_091_module_data_out[4] ,
    \sw_091_module_data_out[3] ,
    \sw_091_module_data_out[2] ,
    \sw_091_module_data_out[1] ,
    \sw_091_module_data_out[0] }));
 user_module_341608574336631379 user_module_341608574336631379_092 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_092_module_data_in[7] ,
    \sw_092_module_data_in[6] ,
    \sw_092_module_data_in[5] ,
    \sw_092_module_data_in[4] ,
    \sw_092_module_data_in[3] ,
    \sw_092_module_data_in[2] ,
    \sw_092_module_data_in[1] ,
    \sw_092_module_data_in[0] }),
    .io_out({\sw_092_module_data_out[7] ,
    \sw_092_module_data_out[6] ,
    \sw_092_module_data_out[5] ,
    \sw_092_module_data_out[4] ,
    \sw_092_module_data_out[3] ,
    \sw_092_module_data_out[2] ,
    \sw_092_module_data_out[1] ,
    \sw_092_module_data_out[0] }));
 user_module_341609034095264340 user_module_341609034095264340_070 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_070_module_data_in[7] ,
    \sw_070_module_data_in[6] ,
    \sw_070_module_data_in[5] ,
    \sw_070_module_data_in[4] ,
    \sw_070_module_data_in[3] ,
    \sw_070_module_data_in[2] ,
    \sw_070_module_data_in[1] ,
    \sw_070_module_data_in[0] }),
    .io_out({\sw_070_module_data_out[7] ,
    \sw_070_module_data_out[6] ,
    \sw_070_module_data_out[5] ,
    \sw_070_module_data_out[4] ,
    \sw_070_module_data_out[3] ,
    \sw_070_module_data_out[2] ,
    \sw_070_module_data_out[1] ,
    \sw_070_module_data_out[0] }));
 user_module_341613097060926036 user_module_341613097060926036_153 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_153_module_data_in[7] ,
    \sw_153_module_data_in[6] ,
    \sw_153_module_data_in[5] ,
    \sw_153_module_data_in[4] ,
    \sw_153_module_data_in[3] ,
    \sw_153_module_data_in[2] ,
    \sw_153_module_data_in[1] ,
    \sw_153_module_data_in[0] }),
    .io_out({\sw_153_module_data_out[7] ,
    \sw_153_module_data_out[6] ,
    \sw_153_module_data_out[5] ,
    \sw_153_module_data_out[4] ,
    \sw_153_module_data_out[3] ,
    \sw_153_module_data_out[2] ,
    \sw_153_module_data_out[1] ,
    \sw_153_module_data_out[0] }));
 user_module_341614346808328788 user_module_341614346808328788_111 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_111_module_data_in[7] ,
    \sw_111_module_data_in[6] ,
    \sw_111_module_data_in[5] ,
    \sw_111_module_data_in[4] ,
    \sw_111_module_data_in[3] ,
    \sw_111_module_data_in[2] ,
    \sw_111_module_data_in[1] ,
    \sw_111_module_data_in[0] }),
    .io_out({\sw_111_module_data_out[7] ,
    \sw_111_module_data_out[6] ,
    \sw_111_module_data_out[5] ,
    \sw_111_module_data_out[4] ,
    \sw_111_module_data_out[3] ,
    \sw_111_module_data_out[2] ,
    \sw_111_module_data_out[1] ,
    \sw_111_module_data_out[0] }));
 user_module_341614374571475540 user_module_341614374571475540_044 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_044_module_data_in[7] ,
    \sw_044_module_data_in[6] ,
    \sw_044_module_data_in[5] ,
    \sw_044_module_data_in[4] ,
    \sw_044_module_data_in[3] ,
    \sw_044_module_data_in[2] ,
    \sw_044_module_data_in[1] ,
    \sw_044_module_data_in[0] }),
    .io_out({\sw_044_module_data_out[7] ,
    \sw_044_module_data_out[6] ,
    \sw_044_module_data_out[5] ,
    \sw_044_module_data_out[4] ,
    \sw_044_module_data_out[3] ,
    \sw_044_module_data_out[2] ,
    \sw_044_module_data_out[1] ,
    \sw_044_module_data_out[0] }));
 user_module_341620484740219475 user_module_341620484740219475_041 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_041_module_data_in[7] ,
    \sw_041_module_data_in[6] ,
    \sw_041_module_data_in[5] ,
    \sw_041_module_data_in[4] ,
    \sw_041_module_data_in[3] ,
    \sw_041_module_data_in[2] ,
    \sw_041_module_data_in[1] ,
    \sw_041_module_data_in[0] }),
    .io_out({\sw_041_module_data_out[7] ,
    \sw_041_module_data_out[6] ,
    \sw_041_module_data_out[5] ,
    \sw_041_module_data_out[4] ,
    \sw_041_module_data_out[3] ,
    \sw_041_module_data_out[2] ,
    \sw_041_module_data_out[1] ,
    \sw_041_module_data_out[0] }));
 user_module_341628725785264722 user_module_341628725785264722_132 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_132_module_data_in[7] ,
    \sw_132_module_data_in[6] ,
    \sw_132_module_data_in[5] ,
    \sw_132_module_data_in[4] ,
    \sw_132_module_data_in[3] ,
    \sw_132_module_data_in[2] ,
    \sw_132_module_data_in[1] ,
    \sw_132_module_data_in[0] }),
    .io_out({\sw_132_module_data_out[7] ,
    \sw_132_module_data_out[6] ,
    \sw_132_module_data_out[5] ,
    \sw_132_module_data_out[4] ,
    \sw_132_module_data_out[3] ,
    \sw_132_module_data_out[2] ,
    \sw_132_module_data_out[1] ,
    \sw_132_module_data_out[0] }));
 user_module_341631511790879314 user_module_341631511790879314_112 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_112_module_data_in[7] ,
    \sw_112_module_data_in[6] ,
    \sw_112_module_data_in[5] ,
    \sw_112_module_data_in[4] ,
    \sw_112_module_data_in[3] ,
    \sw_112_module_data_in[2] ,
    \sw_112_module_data_in[1] ,
    \sw_112_module_data_in[0] }),
    .io_out({\sw_112_module_data_out[7] ,
    \sw_112_module_data_out[6] ,
    \sw_112_module_data_out[5] ,
    \sw_112_module_data_out[4] ,
    \sw_112_module_data_out[3] ,
    \sw_112_module_data_out[2] ,
    \sw_112_module_data_out[1] ,
    \sw_112_module_data_out[0] }));
 user_module_341631644820570706 user_module_341631644820570706_136 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_136_module_data_in[7] ,
    \sw_136_module_data_in[6] ,
    \sw_136_module_data_in[5] ,
    \sw_136_module_data_in[4] ,
    \sw_136_module_data_in[3] ,
    \sw_136_module_data_in[2] ,
    \sw_136_module_data_in[1] ,
    \sw_136_module_data_in[0] }),
    .io_out({\sw_136_module_data_out[7] ,
    \sw_136_module_data_out[6] ,
    \sw_136_module_data_out[5] ,
    \sw_136_module_data_out[4] ,
    \sw_136_module_data_out[3] ,
    \sw_136_module_data_out[2] ,
    \sw_136_module_data_out[1] ,
    \sw_136_module_data_out[0] }));
 user_module_341678527574180436 user_module_341678527574180436_158 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_158_module_data_in[7] ,
    \sw_158_module_data_in[6] ,
    \sw_158_module_data_in[5] ,
    \sw_158_module_data_in[4] ,
    \sw_158_module_data_in[3] ,
    \sw_158_module_data_in[2] ,
    \sw_158_module_data_in[1] ,
    \sw_158_module_data_in[0] }),
    .io_out({\sw_158_module_data_out[7] ,
    \sw_158_module_data_out[6] ,
    \sw_158_module_data_out[5] ,
    \sw_158_module_data_out[4] ,
    \sw_158_module_data_out[3] ,
    \sw_158_module_data_out[2] ,
    \sw_158_module_data_out[1] ,
    \sw_158_module_data_out[0] }));
 user_module_342981109408072274 user_module_342981109408072274_022 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_022_module_data_in[7] ,
    \sw_022_module_data_in[6] ,
    \sw_022_module_data_in[5] ,
    \sw_022_module_data_in[4] ,
    \sw_022_module_data_in[3] ,
    \sw_022_module_data_in[2] ,
    \sw_022_module_data_in[1] ,
    \sw_022_module_data_in[0] }),
    .io_out({\sw_022_module_data_out[7] ,
    \sw_022_module_data_out[6] ,
    \sw_022_module_data_out[5] ,
    \sw_022_module_data_out[4] ,
    \sw_022_module_data_out[3] ,
    \sw_022_module_data_out[2] ,
    \sw_022_module_data_out[1] ,
    \sw_022_module_data_out[0] }));
 user_module_346553315158393428 user_module_346553315158393428_016 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_016_module_data_in[7] ,
    \sw_016_module_data_in[6] ,
    \sw_016_module_data_in[5] ,
    \sw_016_module_data_in[4] ,
    \sw_016_module_data_in[3] ,
    \sw_016_module_data_in[2] ,
    \sw_016_module_data_in[1] ,
    \sw_016_module_data_in[0] }),
    .io_out({\sw_016_module_data_out[7] ,
    \sw_016_module_data_out[6] ,
    \sw_016_module_data_out[5] ,
    \sw_016_module_data_out[4] ,
    \sw_016_module_data_out[3] ,
    \sw_016_module_data_out[2] ,
    \sw_016_module_data_out[1] ,
    \sw_016_module_data_out[0] }));
 user_module_346916357828248146 user_module_346916357828248146_018 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_018_module_data_in[7] ,
    \sw_018_module_data_in[6] ,
    \sw_018_module_data_in[5] ,
    \sw_018_module_data_in[4] ,
    \sw_018_module_data_in[3] ,
    \sw_018_module_data_in[2] ,
    \sw_018_module_data_in[1] ,
    \sw_018_module_data_in[0] }),
    .io_out({\sw_018_module_data_out[7] ,
    \sw_018_module_data_out[6] ,
    \sw_018_module_data_out[5] ,
    \sw_018_module_data_out[4] ,
    \sw_018_module_data_out[3] ,
    \sw_018_module_data_out[2] ,
    \sw_018_module_data_out[1] ,
    \sw_018_module_data_out[0] }));
 user_module_347140425276981843 user_module_347140425276981843_161 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_161_module_data_in[7] ,
    \sw_161_module_data_in[6] ,
    \sw_161_module_data_in[5] ,
    \sw_161_module_data_in[4] ,
    \sw_161_module_data_in[3] ,
    \sw_161_module_data_in[2] ,
    \sw_161_module_data_in[1] ,
    \sw_161_module_data_in[0] }),
    .io_out({\sw_161_module_data_out[7] ,
    \sw_161_module_data_out[6] ,
    \sw_161_module_data_out[5] ,
    \sw_161_module_data_out[4] ,
    \sw_161_module_data_out[3] ,
    \sw_161_module_data_out[2] ,
    \sw_161_module_data_out[1] ,
    \sw_161_module_data_out[0] }));
 user_module_347144898258928211 user_module_347144898258928211_162 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_162_module_data_in[7] ,
    \sw_162_module_data_in[6] ,
    \sw_162_module_data_in[5] ,
    \sw_162_module_data_in[4] ,
    \sw_162_module_data_in[3] ,
    \sw_162_module_data_in[2] ,
    \sw_162_module_data_in[1] ,
    \sw_162_module_data_in[0] }),
    .io_out({\sw_162_module_data_out[7] ,
    \sw_162_module_data_out[6] ,
    \sw_162_module_data_out[5] ,
    \sw_162_module_data_out[4] ,
    \sw_162_module_data_out[3] ,
    \sw_162_module_data_out[2] ,
    \sw_162_module_data_out[1] ,
    \sw_162_module_data_out[0] }));
 user_module_347417602591556180 user_module_347417602591556180_163 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_163_module_data_in[7] ,
    \sw_163_module_data_in[6] ,
    \sw_163_module_data_in[5] ,
    \sw_163_module_data_in[4] ,
    \sw_163_module_data_in[3] ,
    \sw_163_module_data_in[2] ,
    \sw_163_module_data_in[1] ,
    \sw_163_module_data_in[0] }),
    .io_out({\sw_163_module_data_out[7] ,
    \sw_163_module_data_out[6] ,
    \sw_163_module_data_out[5] ,
    \sw_163_module_data_out[4] ,
    \sw_163_module_data_out[3] ,
    \sw_163_module_data_out[2] ,
    \sw_163_module_data_out[1] ,
    \sw_163_module_data_out[0] }));
 user_module_347497504164545108 user_module_347497504164545108_160 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_160_module_data_in[7] ,
    \sw_160_module_data_in[6] ,
    \sw_160_module_data_in[5] ,
    \sw_160_module_data_in[4] ,
    \sw_160_module_data_in[3] ,
    \sw_160_module_data_in[2] ,
    \sw_160_module_data_in[1] ,
    \sw_160_module_data_in[0] }),
    .io_out({\sw_160_module_data_out[7] ,
    \sw_160_module_data_out[6] ,
    \sw_160_module_data_out[5] ,
    \sw_160_module_data_out[4] ,
    \sw_160_module_data_out[3] ,
    \sw_160_module_data_out[2] ,
    \sw_160_module_data_out[1] ,
    \sw_160_module_data_out[0] }));
 user_module_347592305412145748 user_module_347592305412145748_013 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_013_module_data_in[7] ,
    \sw_013_module_data_in[6] ,
    \sw_013_module_data_in[5] ,
    \sw_013_module_data_in[4] ,
    \sw_013_module_data_in[3] ,
    \sw_013_module_data_in[2] ,
    \sw_013_module_data_in[1] ,
    \sw_013_module_data_in[0] }),
    .io_out({\sw_013_module_data_out[7] ,
    \sw_013_module_data_out[6] ,
    \sw_013_module_data_out[5] ,
    \sw_013_module_data_out[4] ,
    \sw_013_module_data_out[3] ,
    \sw_013_module_data_out[2] ,
    \sw_013_module_data_out[1] ,
    \sw_013_module_data_out[0] }));
 user_module_347594509754827347 user_module_347594509754827347_019 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_019_module_data_in[7] ,
    \sw_019_module_data_in[6] ,
    \sw_019_module_data_in[5] ,
    \sw_019_module_data_in[4] ,
    \sw_019_module_data_in[3] ,
    \sw_019_module_data_in[2] ,
    \sw_019_module_data_in[1] ,
    \sw_019_module_data_in[0] }),
    .io_out({\sw_019_module_data_out[7] ,
    \sw_019_module_data_out[6] ,
    \sw_019_module_data_out[5] ,
    \sw_019_module_data_out[4] ,
    \sw_019_module_data_out[3] ,
    \sw_019_module_data_out[2] ,
    \sw_019_module_data_out[1] ,
    \sw_019_module_data_out[0] }));
 user_module_347619669052490324 user_module_347619669052490324_057 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_057_module_data_in[7] ,
    \sw_057_module_data_in[6] ,
    \sw_057_module_data_in[5] ,
    \sw_057_module_data_in[4] ,
    \sw_057_module_data_in[3] ,
    \sw_057_module_data_in[2] ,
    \sw_057_module_data_in[1] ,
    \sw_057_module_data_in[0] }),
    .io_out({\sw_057_module_data_out[7] ,
    \sw_057_module_data_out[6] ,
    \sw_057_module_data_out[5] ,
    \sw_057_module_data_out[4] ,
    \sw_057_module_data_out[3] ,
    \sw_057_module_data_out[2] ,
    \sw_057_module_data_out[1] ,
    \sw_057_module_data_out[0] }));
 user_module_347688030570545747 user_module_347688030570545747_021 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_021_module_data_in[7] ,
    \sw_021_module_data_in[6] ,
    \sw_021_module_data_in[5] ,
    \sw_021_module_data_in[4] ,
    \sw_021_module_data_in[3] ,
    \sw_021_module_data_in[2] ,
    \sw_021_module_data_in[1] ,
    \sw_021_module_data_in[0] }),
    .io_out({\sw_021_module_data_out[7] ,
    \sw_021_module_data_out[6] ,
    \sw_021_module_data_out[5] ,
    \sw_021_module_data_out[4] ,
    \sw_021_module_data_out[3] ,
    \sw_021_module_data_out[2] ,
    \sw_021_module_data_out[1] ,
    \sw_021_module_data_out[0] }));
 user_module_347690870424732244 user_module_347690870424732244_012 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_012_module_data_in[7] ,
    \sw_012_module_data_in[6] ,
    \sw_012_module_data_in[5] ,
    \sw_012_module_data_in[4] ,
    \sw_012_module_data_in[3] ,
    \sw_012_module_data_in[2] ,
    \sw_012_module_data_in[1] ,
    \sw_012_module_data_in[0] }),
    .io_out({\sw_012_module_data_out[7] ,
    \sw_012_module_data_out[6] ,
    \sw_012_module_data_out[5] ,
    \sw_012_module_data_out[4] ,
    \sw_012_module_data_out[3] ,
    \sw_012_module_data_out[2] ,
    \sw_012_module_data_out[1] ,
    \sw_012_module_data_out[0] }));
 user_module_347787021138264660 user_module_347787021138264660_010 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_010_module_data_in[7] ,
    \sw_010_module_data_in[6] ,
    \sw_010_module_data_in[5] ,
    \sw_010_module_data_in[4] ,
    \sw_010_module_data_in[3] ,
    \sw_010_module_data_in[2] ,
    \sw_010_module_data_in[1] ,
    \sw_010_module_data_in[0] }),
    .io_out({\sw_010_module_data_out[7] ,
    \sw_010_module_data_out[6] ,
    \sw_010_module_data_out[5] ,
    \sw_010_module_data_out[4] ,
    \sw_010_module_data_out[3] ,
    \sw_010_module_data_out[2] ,
    \sw_010_module_data_out[1] ,
    \sw_010_module_data_out[0] }));
 user_module_347894637149553236 user_module_347894637149553236_017 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_017_module_data_in[7] ,
    \sw_017_module_data_in[6] ,
    \sw_017_module_data_in[5] ,
    \sw_017_module_data_in[4] ,
    \sw_017_module_data_in[3] ,
    \sw_017_module_data_in[2] ,
    \sw_017_module_data_in[1] ,
    \sw_017_module_data_in[0] }),
    .io_out({\sw_017_module_data_out[7] ,
    \sw_017_module_data_out[6] ,
    \sw_017_module_data_out[5] ,
    \sw_017_module_data_out[4] ,
    \sw_017_module_data_out[3] ,
    \sw_017_module_data_out[2] ,
    \sw_017_module_data_out[1] ,
    \sw_017_module_data_out[0] }));
 user_module_348121131386929746 user_module_348121131386929746_028 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_028_module_data_in[7] ,
    \sw_028_module_data_in[6] ,
    \sw_028_module_data_in[5] ,
    \sw_028_module_data_in[4] ,
    \sw_028_module_data_in[3] ,
    \sw_028_module_data_in[2] ,
    \sw_028_module_data_in[1] ,
    \sw_028_module_data_in[0] }),
    .io_out({\sw_028_module_data_out[7] ,
    \sw_028_module_data_out[6] ,
    \sw_028_module_data_out[5] ,
    \sw_028_module_data_out[4] ,
    \sw_028_module_data_out[3] ,
    \sw_028_module_data_out[2] ,
    \sw_028_module_data_out[1] ,
    \sw_028_module_data_out[0] }));
 user_module_348195845106041428 user_module_348195845106041428_027 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_027_module_data_in[7] ,
    \sw_027_module_data_in[6] ,
    \sw_027_module_data_in[5] ,
    \sw_027_module_data_in[4] ,
    \sw_027_module_data_in[3] ,
    \sw_027_module_data_in[2] ,
    \sw_027_module_data_in[1] ,
    \sw_027_module_data_in[0] }),
    .io_out({\sw_027_module_data_out[7] ,
    \sw_027_module_data_out[6] ,
    \sw_027_module_data_out[5] ,
    \sw_027_module_data_out[4] ,
    \sw_027_module_data_out[3] ,
    \sw_027_module_data_out[2] ,
    \sw_027_module_data_out[1] ,
    \sw_027_module_data_out[0] }));
 user_module_348242239268323922 user_module_348242239268323922_037 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_037_module_data_in[7] ,
    \sw_037_module_data_in[6] ,
    \sw_037_module_data_in[5] ,
    \sw_037_module_data_in[4] ,
    \sw_037_module_data_in[3] ,
    \sw_037_module_data_in[2] ,
    \sw_037_module_data_in[1] ,
    \sw_037_module_data_in[0] }),
    .io_out({\sw_037_module_data_out[7] ,
    \sw_037_module_data_out[6] ,
    \sw_037_module_data_out[5] ,
    \sw_037_module_data_out[4] ,
    \sw_037_module_data_out[3] ,
    \sw_037_module_data_out[2] ,
    \sw_037_module_data_out[1] ,
    \sw_037_module_data_out[0] }));
 user_module_348255968419643987 user_module_348255968419643987_032 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_032_module_data_in[7] ,
    \sw_032_module_data_in[6] ,
    \sw_032_module_data_in[5] ,
    \sw_032_module_data_in[4] ,
    \sw_032_module_data_in[3] ,
    \sw_032_module_data_in[2] ,
    \sw_032_module_data_in[1] ,
    \sw_032_module_data_in[0] }),
    .io_out({\sw_032_module_data_out[7] ,
    \sw_032_module_data_out[6] ,
    \sw_032_module_data_out[5] ,
    \sw_032_module_data_out[4] ,
    \sw_032_module_data_out[3] ,
    \sw_032_module_data_out[2] ,
    \sw_032_module_data_out[1] ,
    \sw_032_module_data_out[0] }));
 user_module_348260124451668562 user_module_348260124451668562_034 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_034_module_data_in[7] ,
    \sw_034_module_data_in[6] ,
    \sw_034_module_data_in[5] ,
    \sw_034_module_data_in[4] ,
    \sw_034_module_data_in[3] ,
    \sw_034_module_data_in[2] ,
    \sw_034_module_data_in[1] ,
    \sw_034_module_data_in[0] }),
    .io_out({\sw_034_module_data_out[7] ,
    \sw_034_module_data_out[6] ,
    \sw_034_module_data_out[5] ,
    \sw_034_module_data_out[4] ,
    \sw_034_module_data_out[3] ,
    \sw_034_module_data_out[2] ,
    \sw_034_module_data_out[1] ,
    \sw_034_module_data_out[0] }));
 user_module_348381622440034899 user_module_348381622440034899_084 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_084_module_data_in[7] ,
    \sw_084_module_data_in[6] ,
    \sw_084_module_data_in[5] ,
    \sw_084_module_data_in[4] ,
    \sw_084_module_data_in[3] ,
    \sw_084_module_data_in[2] ,
    \sw_084_module_data_in[1] ,
    \sw_084_module_data_in[0] }),
    .io_out({\sw_084_module_data_out[7] ,
    \sw_084_module_data_out[6] ,
    \sw_084_module_data_out[5] ,
    \sw_084_module_data_out[4] ,
    \sw_084_module_data_out[3] ,
    \sw_084_module_data_out[2] ,
    \sw_084_module_data_out[1] ,
    \sw_084_module_data_out[0] }));
 user_module_348540666182107731 user_module_348540666182107731_064 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_064_module_data_in[7] ,
    \sw_064_module_data_in[6] ,
    \sw_064_module_data_in[5] ,
    \sw_064_module_data_in[4] ,
    \sw_064_module_data_in[3] ,
    \sw_064_module_data_in[2] ,
    \sw_064_module_data_in[1] ,
    \sw_064_module_data_in[0] }),
    .io_out({\sw_064_module_data_out[7] ,
    \sw_064_module_data_out[6] ,
    \sw_064_module_data_out[5] ,
    \sw_064_module_data_out[4] ,
    \sw_064_module_data_out[3] ,
    \sw_064_module_data_out[2] ,
    \sw_064_module_data_out[1] ,
    \sw_064_module_data_out[0] }));
 user_module_348787952842703444 user_module_348787952842703444_096 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_096_module_data_in[7] ,
    \sw_096_module_data_in[6] ,
    \sw_096_module_data_in[5] ,
    \sw_096_module_data_in[4] ,
    \sw_096_module_data_in[3] ,
    \sw_096_module_data_in[2] ,
    \sw_096_module_data_in[1] ,
    \sw_096_module_data_in[0] }),
    .io_out({\sw_096_module_data_out[7] ,
    \sw_096_module_data_out[6] ,
    \sw_096_module_data_out[5] ,
    \sw_096_module_data_out[4] ,
    \sw_096_module_data_out[3] ,
    \sw_096_module_data_out[2] ,
    \sw_096_module_data_out[1] ,
    \sw_096_module_data_out[0] }));
 user_module_349011320806310484 user_module_349011320806310484_072 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_072_module_data_in[7] ,
    \sw_072_module_data_in[6] ,
    \sw_072_module_data_in[5] ,
    \sw_072_module_data_in[4] ,
    \sw_072_module_data_in[3] ,
    \sw_072_module_data_in[2] ,
    \sw_072_module_data_in[1] ,
    \sw_072_module_data_in[0] }),
    .io_out({\sw_072_module_data_out[7] ,
    \sw_072_module_data_out[6] ,
    \sw_072_module_data_out[5] ,
    \sw_072_module_data_out[4] ,
    \sw_072_module_data_out[3] ,
    \sw_072_module_data_out[2] ,
    \sw_072_module_data_out[1] ,
    \sw_072_module_data_out[0] }));
 user_module_349047610915422802 user_module_349047610915422802_066 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_066_module_data_in[7] ,
    \sw_066_module_data_in[6] ,
    \sw_066_module_data_in[5] ,
    \sw_066_module_data_in[4] ,
    \sw_066_module_data_in[3] ,
    \sw_066_module_data_in[2] ,
    \sw_066_module_data_in[1] ,
    \sw_066_module_data_in[0] }),
    .io_out({\sw_066_module_data_out[7] ,
    \sw_066_module_data_out[6] ,
    \sw_066_module_data_out[5] ,
    \sw_066_module_data_out[4] ,
    \sw_066_module_data_out[3] ,
    \sw_066_module_data_out[2] ,
    \sw_066_module_data_out[1] ,
    \sw_066_module_data_out[0] }));
 user_module_349228308755382868 user_module_349228308755382868_082 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_082_module_data_in[7] ,
    \sw_082_module_data_in[6] ,
    \sw_082_module_data_in[5] ,
    \sw_082_module_data_in[4] ,
    \sw_082_module_data_in[3] ,
    \sw_082_module_data_in[2] ,
    \sw_082_module_data_in[1] ,
    \sw_082_module_data_in[0] }),
    .io_out({\sw_082_module_data_out[7] ,
    \sw_082_module_data_out[6] ,
    \sw_082_module_data_out[5] ,
    \sw_082_module_data_out[4] ,
    \sw_082_module_data_out[3] ,
    \sw_082_module_data_out[2] ,
    \sw_082_module_data_out[1] ,
    \sw_082_module_data_out[0] }));
 user_module_349255310782759507 user_module_349255310782759507_126 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_126_module_data_in[7] ,
    \sw_126_module_data_in[6] ,
    \sw_126_module_data_in[5] ,
    \sw_126_module_data_in[4] ,
    \sw_126_module_data_in[3] ,
    \sw_126_module_data_in[2] ,
    \sw_126_module_data_in[1] ,
    \sw_126_module_data_in[0] }),
    .io_out({\sw_126_module_data_out[7] ,
    \sw_126_module_data_out[6] ,
    \sw_126_module_data_out[5] ,
    \sw_126_module_data_out[4] ,
    \sw_126_module_data_out[3] ,
    \sw_126_module_data_out[2] ,
    \sw_126_module_data_out[1] ,
    \sw_126_module_data_out[0] }));
 user_module_349519263900369490 user_module_349519263900369490_146 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_146_module_data_in[7] ,
    \sw_146_module_data_in[6] ,
    \sw_146_module_data_in[5] ,
    \sw_146_module_data_in[4] ,
    \sw_146_module_data_in[3] ,
    \sw_146_module_data_in[2] ,
    \sw_146_module_data_in[1] ,
    \sw_146_module_data_in[0] }),
    .io_out({\sw_146_module_data_out[7] ,
    \sw_146_module_data_out[6] ,
    \sw_146_module_data_out[5] ,
    \sw_146_module_data_out[4] ,
    \sw_146_module_data_out[3] ,
    \sw_146_module_data_out[2] ,
    \sw_146_module_data_out[1] ,
    \sw_146_module_data_out[0] }));
 user_module_349546262775726676 user_module_349546262775726676_087 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_087_module_data_in[7] ,
    \sw_087_module_data_in[6] ,
    \sw_087_module_data_in[5] ,
    \sw_087_module_data_in[4] ,
    \sw_087_module_data_in[3] ,
    \sw_087_module_data_in[2] ,
    \sw_087_module_data_in[1] ,
    \sw_087_module_data_in[0] }),
    .io_out({\sw_087_module_data_out[7] ,
    \sw_087_module_data_out[6] ,
    \sw_087_module_data_out[5] ,
    \sw_087_module_data_out[4] ,
    \sw_087_module_data_out[3] ,
    \sw_087_module_data_out[2] ,
    \sw_087_module_data_out[1] ,
    \sw_087_module_data_out[0] }));
 user_module_349729432862196307 user_module_349729432862196307_105 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_105_module_data_in[7] ,
    \sw_105_module_data_in[6] ,
    \sw_105_module_data_in[5] ,
    \sw_105_module_data_in[4] ,
    \sw_105_module_data_in[3] ,
    \sw_105_module_data_in[2] ,
    \sw_105_module_data_in[1] ,
    \sw_105_module_data_in[0] }),
    .io_out({\sw_105_module_data_out[7] ,
    \sw_105_module_data_out[6] ,
    \sw_105_module_data_out[5] ,
    \sw_105_module_data_out[4] ,
    \sw_105_module_data_out[3] ,
    \sw_105_module_data_out[2] ,
    \sw_105_module_data_out[1] ,
    \sw_105_module_data_out[0] }));
 user_module_349790606404354643 user_module_349790606404354643_102 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_102_module_data_in[7] ,
    \sw_102_module_data_in[6] ,
    \sw_102_module_data_in[5] ,
    \sw_102_module_data_in[4] ,
    \sw_102_module_data_in[3] ,
    \sw_102_module_data_in[2] ,
    \sw_102_module_data_in[1] ,
    \sw_102_module_data_in[0] }),
    .io_out({\sw_102_module_data_out[7] ,
    \sw_102_module_data_out[6] ,
    \sw_102_module_data_out[5] ,
    \sw_102_module_data_out[4] ,
    \sw_102_module_data_out[3] ,
    \sw_102_module_data_out[2] ,
    \sw_102_module_data_out[1] ,
    \sw_102_module_data_out[0] }));
 user_module_349803790984020562 user_module_349803790984020562_148 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_148_module_data_in[7] ,
    \sw_148_module_data_in[6] ,
    \sw_148_module_data_in[5] ,
    \sw_148_module_data_in[4] ,
    \sw_148_module_data_in[3] ,
    \sw_148_module_data_in[2] ,
    \sw_148_module_data_in[1] ,
    \sw_148_module_data_in[0] }),
    .io_out({\sw_148_module_data_out[7] ,
    \sw_148_module_data_out[6] ,
    \sw_148_module_data_out[5] ,
    \sw_148_module_data_out[4] ,
    \sw_148_module_data_out[3] ,
    \sw_148_module_data_out[2] ,
    \sw_148_module_data_out[1] ,
    \sw_148_module_data_out[0] }));
 user_module_349813388252021330 user_module_349813388252021330_129 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_129_module_data_in[7] ,
    \sw_129_module_data_in[6] ,
    \sw_129_module_data_in[5] ,
    \sw_129_module_data_in[4] ,
    \sw_129_module_data_in[3] ,
    \sw_129_module_data_in[2] ,
    \sw_129_module_data_in[1] ,
    \sw_129_module_data_in[0] }),
    .io_out({\sw_129_module_data_out[7] ,
    \sw_129_module_data_out[6] ,
    \sw_129_module_data_out[5] ,
    \sw_129_module_data_out[4] ,
    \sw_129_module_data_out[3] ,
    \sw_129_module_data_out[2] ,
    \sw_129_module_data_out[1] ,
    \sw_129_module_data_out[0] }));
 user_module_349833797657690706 user_module_349833797657690706_134 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_134_module_data_in[7] ,
    \sw_134_module_data_in[6] ,
    \sw_134_module_data_in[5] ,
    \sw_134_module_data_in[4] ,
    \sw_134_module_data_in[3] ,
    \sw_134_module_data_in[2] ,
    \sw_134_module_data_in[1] ,
    \sw_134_module_data_in[0] }),
    .io_out({\sw_134_module_data_out[7] ,
    \sw_134_module_data_out[6] ,
    \sw_134_module_data_out[5] ,
    \sw_134_module_data_out[4] ,
    \sw_134_module_data_out[3] ,
    \sw_134_module_data_out[2] ,
    \sw_134_module_data_out[1] ,
    \sw_134_module_data_out[0] }));
 user_module_349886696875098706 user_module_349886696875098706_117 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_117_module_data_in[7] ,
    \sw_117_module_data_in[6] ,
    \sw_117_module_data_in[5] ,
    \sw_117_module_data_in[4] ,
    \sw_117_module_data_in[3] ,
    \sw_117_module_data_in[2] ,
    \sw_117_module_data_in[1] ,
    \sw_117_module_data_in[0] }),
    .io_out({\sw_117_module_data_out[7] ,
    \sw_117_module_data_out[6] ,
    \sw_117_module_data_out[5] ,
    \sw_117_module_data_out[4] ,
    \sw_117_module_data_out[3] ,
    \sw_117_module_data_out[2] ,
    \sw_117_module_data_out[1] ,
    \sw_117_module_data_out[0] }));
 user_module_349901899339661908 user_module_349901899339661908_062 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_062_module_data_in[7] ,
    \sw_062_module_data_in[6] ,
    \sw_062_module_data_in[5] ,
    \sw_062_module_data_in[4] ,
    \sw_062_module_data_in[3] ,
    \sw_062_module_data_in[2] ,
    \sw_062_module_data_in[1] ,
    \sw_062_module_data_in[0] }),
    .io_out({\sw_062_module_data_out[7] ,
    \sw_062_module_data_out[6] ,
    \sw_062_module_data_out[5] ,
    \sw_062_module_data_out[4] ,
    \sw_062_module_data_out[3] ,
    \sw_062_module_data_out[2] ,
    \sw_062_module_data_out[1] ,
    \sw_062_module_data_out[0] }));
 user_module_349934460979905106 user_module_349934460979905106_130 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_130_module_data_in[7] ,
    \sw_130_module_data_in[6] ,
    \sw_130_module_data_in[5] ,
    \sw_130_module_data_in[4] ,
    \sw_130_module_data_in[3] ,
    \sw_130_module_data_in[2] ,
    \sw_130_module_data_in[1] ,
    \sw_130_module_data_in[0] }),
    .io_out({\sw_130_module_data_out[7] ,
    \sw_130_module_data_out[6] ,
    \sw_130_module_data_out[5] ,
    \sw_130_module_data_out[4] ,
    \sw_130_module_data_out[3] ,
    \sw_130_module_data_out[2] ,
    \sw_130_module_data_out[1] ,
    \sw_130_module_data_out[0] }));
 user_module_349952820323025491 user_module_349952820323025491_142 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_142_module_data_in[7] ,
    \sw_142_module_data_in[6] ,
    \sw_142_module_data_in[5] ,
    \sw_142_module_data_in[4] ,
    \sw_142_module_data_in[3] ,
    \sw_142_module_data_in[2] ,
    \sw_142_module_data_in[1] ,
    \sw_142_module_data_in[0] }),
    .io_out({\sw_142_module_data_out[7] ,
    \sw_142_module_data_out[6] ,
    \sw_142_module_data_out[5] ,
    \sw_142_module_data_out[4] ,
    \sw_142_module_data_out[3] ,
    \sw_142_module_data_out[2] ,
    \sw_142_module_data_out[1] ,
    \sw_142_module_data_out[0] }));
 user_module_349953952950780498 user_module_349953952950780498_063 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_063_module_data_in[7] ,
    \sw_063_module_data_in[6] ,
    \sw_063_module_data_in[5] ,
    \sw_063_module_data_in[4] ,
    \sw_063_module_data_in[3] ,
    \sw_063_module_data_in[2] ,
    \sw_063_module_data_in[1] ,
    \sw_063_module_data_in[0] }),
    .io_out({\sw_063_module_data_out[7] ,
    \sw_063_module_data_out[6] ,
    \sw_063_module_data_out[5] ,
    \sw_063_module_data_out[4] ,
    \sw_063_module_data_out[3] ,
    \sw_063_module_data_out[2] ,
    \sw_063_module_data_out[1] ,
    \sw_063_module_data_out[0] }));
 user_module_nickoe user_module_nickoe_059 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_059_module_data_in[7] ,
    \sw_059_module_data_in[6] ,
    \sw_059_module_data_in[5] ,
    \sw_059_module_data_in[4] ,
    \sw_059_module_data_in[3] ,
    \sw_059_module_data_in[2] ,
    \sw_059_module_data_in[1] ,
    \sw_059_module_data_in[0] }),
    .io_out({\sw_059_module_data_out[7] ,
    \sw_059_module_data_out[6] ,
    \sw_059_module_data_out[5] ,
    \sw_059_module_data_out[4] ,
    \sw_059_module_data_out[3] ,
    \sw_059_module_data_out[2] ,
    \sw_059_module_data_out[1] ,
    \sw_059_module_data_out[0] }));
 user_module_skylersaleh user_module_skylersaleh_131 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_131_module_data_in[7] ,
    \sw_131_module_data_in[6] ,
    \sw_131_module_data_in[5] ,
    \sw_131_module_data_in[4] ,
    \sw_131_module_data_in[3] ,
    \sw_131_module_data_in[2] ,
    \sw_131_module_data_in[1] ,
    \sw_131_module_data_in[0] }),
    .io_out({\sw_131_module_data_out[7] ,
    \sw_131_module_data_out[6] ,
    \sw_131_module_data_out[5] ,
    \sw_131_module_data_out[4] ,
    \sw_131_module_data_out[3] ,
    \sw_131_module_data_out[2] ,
    \sw_131_module_data_out[1] ,
    \sw_131_module_data_out[0] }));
 vaishnavachath_rotary_toplevel vaishnavachath_rotary_toplevel_110 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_110_module_data_in[7] ,
    \sw_110_module_data_in[6] ,
    \sw_110_module_data_in[5] ,
    \sw_110_module_data_in[4] ,
    \sw_110_module_data_in[3] ,
    \sw_110_module_data_in[2] ,
    \sw_110_module_data_in[1] ,
    \sw_110_module_data_in[0] }),
    .io_out({\sw_110_module_data_out[7] ,
    \sw_110_module_data_out[6] ,
    \sw_110_module_data_out[5] ,
    \sw_110_module_data_out[4] ,
    \sw_110_module_data_out[3] ,
    \sw_110_module_data_out[2] ,
    \sw_110_module_data_out[1] ,
    \sw_110_module_data_out[0] }));
 wren6991_whisk_tt2_io_wrapper wren6991_whisk_tt2_io_wrapper_093 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_093_module_data_in[7] ,
    \sw_093_module_data_in[6] ,
    \sw_093_module_data_in[5] ,
    \sw_093_module_data_in[4] ,
    \sw_093_module_data_in[3] ,
    \sw_093_module_data_in[2] ,
    \sw_093_module_data_in[1] ,
    \sw_093_module_data_in[0] }),
    .io_out({\sw_093_module_data_out[7] ,
    \sw_093_module_data_out[6] ,
    \sw_093_module_data_out[5] ,
    \sw_093_module_data_out[4] ,
    \sw_093_module_data_out[3] ,
    \sw_093_module_data_out[2] ,
    \sw_093_module_data_out[1] ,
    \sw_093_module_data_out[0] }));
 xor_shift32_evango xor_shift32_evango_053 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_053_module_data_in[7] ,
    \sw_053_module_data_in[6] ,
    \sw_053_module_data_in[5] ,
    \sw_053_module_data_in[4] ,
    \sw_053_module_data_in[3] ,
    \sw_053_module_data_in[2] ,
    \sw_053_module_data_in[1] ,
    \sw_053_module_data_in[0] }),
    .io_out({\sw_053_module_data_out[7] ,
    \sw_053_module_data_out[6] ,
    \sw_053_module_data_out[5] ,
    \sw_053_module_data_out[4] ,
    \sw_053_module_data_out[3] ,
    \sw_053_module_data_out[2] ,
    \sw_053_module_data_out[1] ,
    \sw_053_module_data_out[0] }));
 xor_shift32_quantamhd xor_shift32_quantamhd_052 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_052_module_data_in[7] ,
    \sw_052_module_data_in[6] ,
    \sw_052_module_data_in[5] ,
    \sw_052_module_data_in[4] ,
    \sw_052_module_data_in[3] ,
    \sw_052_module_data_in[2] ,
    \sw_052_module_data_in[1] ,
    \sw_052_module_data_in[0] }),
    .io_out({\sw_052_module_data_out[7] ,
    \sw_052_module_data_out[6] ,
    \sw_052_module_data_out[5] ,
    \sw_052_module_data_out[4] ,
    \sw_052_module_data_out[3] ,
    \sw_052_module_data_out[2] ,
    \sw_052_module_data_out[1] ,
    \sw_052_module_data_out[0] }));
 xyz_peppergray_Potato1_top xyz_peppergray_Potato1_top_030 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_030_module_data_in[7] ,
    \sw_030_module_data_in[6] ,
    \sw_030_module_data_in[5] ,
    \sw_030_module_data_in[4] ,
    \sw_030_module_data_in[3] ,
    \sw_030_module_data_in[2] ,
    \sw_030_module_data_in[1] ,
    \sw_030_module_data_in[0] }),
    .io_out({\sw_030_module_data_out[7] ,
    \sw_030_module_data_out[6] ,
    \sw_030_module_data_out[5] ,
    \sw_030_module_data_out[4] ,
    \sw_030_module_data_out[3] ,
    \sw_030_module_data_out[2] ,
    \sw_030_module_data_out[1] ,
    \sw_030_module_data_out[0] }));
 yubex_egg_timer yubex_egg_timer_029 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_029_module_data_in[7] ,
    \sw_029_module_data_in[6] ,
    \sw_029_module_data_in[5] ,
    \sw_029_module_data_in[4] ,
    \sw_029_module_data_in[3] ,
    \sw_029_module_data_in[2] ,
    \sw_029_module_data_in[1] ,
    \sw_029_module_data_in[0] }),
    .io_out({\sw_029_module_data_out[7] ,
    \sw_029_module_data_out[6] ,
    \sw_029_module_data_out[5] ,
    \sw_029_module_data_out[4] ,
    \sw_029_module_data_out[3] ,
    \sw_029_module_data_out[2] ,
    \sw_029_module_data_out[1] ,
    \sw_029_module_data_out[0] }));
 yupferris_bitslam yupferris_bitslam_040 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_040_module_data_in[7] ,
    \sw_040_module_data_in[6] ,
    \sw_040_module_data_in[5] ,
    \sw_040_module_data_in[4] ,
    \sw_040_module_data_in[3] ,
    \sw_040_module_data_in[2] ,
    \sw_040_module_data_in[1] ,
    \sw_040_module_data_in[0] }),
    .io_out({\sw_040_module_data_out[7] ,
    \sw_040_module_data_out[6] ,
    \sw_040_module_data_out[5] ,
    \sw_040_module_data_out[4] ,
    \sw_040_module_data_out[3] ,
    \sw_040_module_data_out[2] ,
    \sw_040_module_data_out[1] ,
    \sw_040_module_data_out[0] }));
 zoechip zoechip_031 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_031_module_data_in[7] ,
    \sw_031_module_data_in[6] ,
    \sw_031_module_data_in[5] ,
    \sw_031_module_data_in[4] ,
    \sw_031_module_data_in[3] ,
    \sw_031_module_data_in[2] ,
    \sw_031_module_data_in[1] ,
    \sw_031_module_data_in[0] }),
    .io_out({\sw_031_module_data_out[7] ,
    \sw_031_module_data_out[6] ,
    \sw_031_module_data_out[5] ,
    \sw_031_module_data_out[4] ,
    \sw_031_module_data_out[3] ,
    \sw_031_module_data_out[2] ,
    \sw_031_module_data_out[1] ,
    \sw_031_module_data_out[0] }));
 zymason_tinytop zymason_tinytop_122 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_122_module_data_in[7] ,
    \sw_122_module_data_in[6] ,
    \sw_122_module_data_in[5] ,
    \sw_122_module_data_in[4] ,
    \sw_122_module_data_in[3] ,
    \sw_122_module_data_in[2] ,
    \sw_122_module_data_in[1] ,
    \sw_122_module_data_in[0] }),
    .io_out({\sw_122_module_data_out[7] ,
    \sw_122_module_data_out[6] ,
    \sw_122_module_data_out[5] ,
    \sw_122_module_data_out[4] ,
    \sw_122_module_data_out[3] ,
    \sw_122_module_data_out[2] ,
    \sw_122_module_data_out[1] ,
    \sw_122_module_data_out[0] }));
endmodule
